`timescale 1ns/1ns

module wt_mem5 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'hfba808fb0668f9cf0d8a066c0826f183e9a5;
mem[1] = 144'h1e00e20c0a96e2f318a60c35facddc4c0fb3;
mem[2] = 144'he52dff27f39b1b79fbe5008a11a2fc8d00a8;
mem[3] = 144'h189fe6510b801a67f0bde8bb12e4f5670e20;
mem[4] = 144'h1ecff7c8f5c0ea6eecaa1cfde6b4ff431ad8;
mem[5] = 144'h0cc2e46409f208d5f45efa18e22b01fa1455;
mem[6] = 144'h0284095c1c7afb050b6aed5f091f08a90d65;
mem[7] = 144'hf6d20bafe13e0ef80d05f52cf910fc38fb2d;
mem[8] = 144'h0566e5350e7defb407f218dc0a9c0a461ed5;
mem[9] = 144'hf325fda81596f2d80964039ef545e194169d;
mem[10] = 144'h0229f5a3e0a9e6fcf2d0e31a14da0fc40abf;
mem[11] = 144'he5dbe730069ff9f112341dbbe6b6f2aafbbf;
mem[12] = 144'h07b9ea50f671e9e110850bcaf86817c0f2d3;
mem[13] = 144'heea30af2fa89e41c0dc5f8bd111c0917141c;
mem[14] = 144'he132021807dc0bc2189ee8b912291993edec;
mem[15] = 144'h19620389eb47e6671167f5a1e2cbf3f2ed75;
mem[16] = 144'h05d10082f6a6f785ff37fc7d13a117b91d64;
mem[17] = 144'he8a1f33af263e0f61be51339039d1ebc1995;
mem[18] = 144'hf4bd18350b07fcf20e01fc620d82e16efc81;
mem[19] = 144'h03460c890efbe9cdfb7cf74003ca15a2fd2d;
mem[20] = 144'h0379ef54fa250b86050fe747f77f177cfc6e;
mem[21] = 144'hfc540228f5c919e70e0bec07e21deb8ef480;
mem[22] = 144'hec2c1bd9e9cdec7df91af98ef5e1f17af7f6;
mem[23] = 144'h05890572ec641ca0f228fc6fe3a814a7f91b;
mem[24] = 144'hf960105802180cec1f441d8703571d18e76c;
mem[25] = 144'hfb8ae5fb1666e2a20638176de2edefb61e08;
mem[26] = 144'h06ea18e416831b2104e8e1ef15970559186f;
mem[27] = 144'hf5d70f2ce17907b4e762fa0d1336146d0e83;
mem[28] = 144'h10631d17f1aef8c8048807c0fb76164d0576;
mem[29] = 144'he71309a7f1ebf397e404180dee55f173fc43;
mem[30] = 144'h02eafc7708340cf9e57f12e71d60e3bf0c31;
mem[31] = 144'h020af5c90509e24b162c1bc114feefb1e2de;
mem[32] = 144'h09c81e73f3321b08ecf9f9a00117e797fb38;
mem[33] = 144'h189e0f461eb3e373fc9cf9b50c76f8effc8c;
mem[34] = 144'hebb611b8072d0f2c002716cf0c96fb450af3;
mem[35] = 144'h01bd05b5fb6e0e6ffbcde0a006f1efa70703;
mem[36] = 144'h127d055ee1840e6cfb06ff9af194e5c1f1f7;
mem[37] = 144'h06f803011597f00b1548ed79e80f15be0332;
mem[38] = 144'h0f200ca1180efcc6044309d90a7907f0178c;
mem[39] = 144'hed450e030051ebf1011e029a15121485ed1f;
mem[40] = 144'h04ac1a961b78eff5188deb4af430129400f7;
mem[41] = 144'h0fd9f8a10e24facaf479fa6b13fa1f2de637;
mem[42] = 144'h09d9f9caef7b14f3189710a3f3b90cd7f292;
mem[43] = 144'he75303e31328f6b4072312e7ef7ef31311f4;
mem[44] = 144'hfc7b0ecafb5016061e3eed3df91801aef4dd;
mem[45] = 144'h11f90b5914e5fdb01e9b0cdbf3db110405f0;
mem[46] = 144'he52710e4fcff03adee7c16810242052d09d2;
mem[47] = 144'h121e0c7bf2d70cf61c4511cbfd91ff7eee7a;
mem[48] = 144'he77216511b2eea5d055204ebf69a0542e0b9;
mem[49] = 144'h0a88f34318fa1d690211fa710a52dff6f37b;
mem[50] = 144'he2a9f844e3541f29002a0e7a0bca10a90ccb;
mem[51] = 144'hefa31f4b17480fec0d8f1a74ec9eeb5a1dd0;
mem[52] = 144'he6ade56bee7c0cb6eda50ceaf944efbd1031;
mem[53] = 144'h0fb1e9a20870e86fff7c0bf9f623138408e4;
mem[54] = 144'hfca7eb2a13eb0d56efb416a61c6d0919f988;
mem[55] = 144'h0d371b661113e06fe07d1faf124214caee6c;
mem[56] = 144'h1111f53800aff218fcfdf863ee6c0f2b19d3;
mem[57] = 144'he75015be1c3df7fc0a65e6f3150b1d5e0957;
mem[58] = 144'h1b320e00e2f0004fe17afafa082004a2fdd3;
mem[59] = 144'h13c01fd31d510d391f0901e61dafe94de4a4;
mem[60] = 144'hfec11a85e62df4690b62001e06611c70e6da;
mem[61] = 144'h01b2edc8064819eee4d0f7c7f9ab1ba40a7d;
mem[62] = 144'hf183f844086e15c6f123f439e487e9ca1d60;
mem[63] = 144'hff6b1e65e9a2f0850e780d1fe25ee97bf870;
mem[64] = 144'h187106b3ffb60f050924f402fa06e8430550;
mem[65] = 144'hea4ee5c6f102081f0275ef730cbf195b163f;
mem[66] = 144'he8380c5704be1f89e84b0abdf905fa7703b5;
mem[67] = 144'h0e9ef71a163b12010b5d143d11ea10c50429;
mem[68] = 144'he7a00dc51e4a09b70c00f3a50741fb93f517;
mem[69] = 144'h1fa60b70e9781b86e60b1d87ffbce117e3da;
mem[70] = 144'he4bcf8ff0bb8038dfadeff1f0cade18b05d5;
mem[71] = 144'hee1a1b9af37e1c96144ff693119a154e1f64;
mem[72] = 144'hf4b811da0c6e129eede20f020707ee990dee;
mem[73] = 144'h1014f716eb9defa2e61119a40bd4111bee7e;
mem[74] = 144'h10b315c913ffec61f1f9e1f8f2e60826e2b3;
mem[75] = 144'hfbdae33d1d440565f748e6e7f9ae01ad1674;
mem[76] = 144'hf1bdfe3f00e5f7c6fbbfff7fe146f4baf2cf;
mem[77] = 144'h03e9e9f0fae410de1f111b5310cef9050d4f;
mem[78] = 144'hf6a4fe9aeabe124d1c7000a1119aeb3cf0b6;
mem[79] = 144'hfebd014e032ced5d02e4f8e61857e681f7ef;
mem[80] = 144'hf747f70c1089efcce9c41eddf521019cefad;
mem[81] = 144'he0ed00e3e66df6201897f916e9afe7f6f12d;
mem[82] = 144'h08c7f932fdd9f8f7ee9a0ee0ee4a1a8cfabb;
mem[83] = 144'hfa94f205fe0f0276e11c022508431bcce469;
mem[84] = 144'hfb95f71ef23307380a82e1b31b601cd00ddb;
mem[85] = 144'he0defde0ea5111e4e1e2e9dbe64d003be5d8;
mem[86] = 144'h154efc4bfd2106b40a31059615c817cde304;
mem[87] = 144'hf83c0b0a1ce20ec5eb40ed6fe8fa10f1f463;
mem[88] = 144'heccf18b6f8f0f437fc4a109a0cc500a40ee8;
mem[89] = 144'h1b87ea34fb7ef627ef8414caed75046bea89;
mem[90] = 144'hf075f1a5fe41030c0439f6bd0351ed3e13a5;
mem[91] = 144'hf21518eaf68210faf3540b4c058be521e72f;
mem[92] = 144'hf941e310e51be260eafbe3691829e3231eb3;
mem[93] = 144'he443e6da18bcf18fecca177308260708f2e4;
mem[94] = 144'hffce18fc115b1ff3103fe67b0d691636e0cb;
mem[95] = 144'h1ab1f5e2e935e8b605250e9cf628ff7d0c75;
mem[96] = 144'hfa8ae85519a2e3d3e37c0debee5b0ccbf4ed;
mem[97] = 144'hfc4b1d71e02c03d0f63be58600501bbfeef6;
mem[98] = 144'h0fc7e831f7f014eaeb960865e868fe8ae71b;
mem[99] = 144'he79802c7f7b4e606ee8303e4e48512e4ea7d;
mem[100] = 144'he94d02f9027c17ec00ac0d781b67e568e203;
mem[101] = 144'hfd2b0da7f091f47c00d00f46f0e7e82d1c73;
mem[102] = 144'hf0400679e56812bbfae6f409f80219fce034;
mem[103] = 144'h08641bb902a4f3f6e1d30ae0e1bcf2e9eb07;
mem[104] = 144'hf60c0a10fb5ff26f083ee4460718e96bf438;
mem[105] = 144'h1eebf6161e71fc890d53fc03ec25e3bcfdc6;
mem[106] = 144'h0bdbe2b7082d1318fcd8041d1ad1116e0b81;
mem[107] = 144'h12f51f2af14901f7fbf3fc8d1241eecb13da;
mem[108] = 144'hef30033f1972ef1c048ef91f115e11fffc3d;
mem[109] = 144'h1c44144700720873e88e12ec190dee6e0ed6;
mem[110] = 144'hf2b7e8c4e007084113861c0618e4fc4e0789;
mem[111] = 144'hfb43f2511a2c0fb319c8ea3401a3e27cea5c;
mem[112] = 144'h00f10b7d02adf1d7f9a5e828fab314e6e125;
mem[113] = 144'hf30c04eb11281ee40ef3fa49eaa31179edb8;
mem[114] = 144'h13890903104b1d180b35fdf9eb281a900366;
mem[115] = 144'h0629fa10e4d718b51a86f62c0a10fd1200ae;
mem[116] = 144'he65ef6e7e0ce12bbfbd215fe1fdbe10def8b;
mem[117] = 144'h0166f299fef606de00ad210dfd3ff45905f1;
mem[118] = 144'heae31f4a1f64e1751c8ef6300218f45804e3;
mem[119] = 144'h0c410ec1e8feea111cd209e70451117012af;
mem[120] = 144'h1190e823ee33f842ef8112f20f86e5aa0aea;
mem[121] = 144'he36ae3030b23e81613ace67e097f1349f624;
mem[122] = 144'h0871fcba04b7f79a167ffe6b0820f5aafe4c;
mem[123] = 144'he85cf7621d550c0ffcbcf7951facfde40ecd;
mem[124] = 144'h1130e46308cafbc81e5318aa163e0e23e9fd;
mem[125] = 144'h00b602eb02961f860572fe2115911f26f096;
mem[126] = 144'h1e021f32f53efb7be78d13881b4013f6f778;
mem[127] = 144'h1bf0122f16eae199eca4fd55efcaeafaee65;
mem[128] = 144'h003108cae98be5b1fe9a187b1cd1052df9ce;
mem[129] = 144'h080bf0ebef76133a1fe8f0910c3413a11cea;
mem[130] = 144'hf14fffe4fd3a193af4d9f4311c0f0009e758;
mem[131] = 144'he0571ae9eae6f07e113203460149f60e02ab;
mem[132] = 144'h00e01c39ea0f0e5df88de331f12c0756f39e;
mem[133] = 144'h1844e2e1fc02e90f12cbfe2e0195f07016be;
mem[134] = 144'hfe93e4d0e2851f670d9a1edb101710b8f66f;
mem[135] = 144'hf6b706431a7e1f60f9041ca90cceed75e365;
mem[136] = 144'h1819e0a8102df6f9e58ae64a0a8c004de753;
mem[137] = 144'h1610f4630f92017c0e70f9b7e868fefc1121;
mem[138] = 144'h02b01ec5029efeade2640175e7c21fecee42;
mem[139] = 144'hf01f09bf18b2021af65ee9f5eded189cea18;
mem[140] = 144'he56ef7da12ff1f4ef6bc078a1d1913321c16;
mem[141] = 144'h1178faf6eadc0482e4351c38f156f2b41a30;
mem[142] = 144'h1234109e161e1b630df1e34af8fef725f9bc;
mem[143] = 144'hf4851e95f2610b0cebde0a47fd7b11a1e66c;
mem[144] = 144'h0ab617fb1625e212ed1bffc9ede7ef32f01c;
mem[145] = 144'hf5ba19f6eae00972e624ec540f4fe8b9126b;
mem[146] = 144'hfbc6e4180d3015d31299090ee2351b5def1b;
mem[147] = 144'h1c20f6d70b01fdaa0222e15a1ca4e88100a4;
mem[148] = 144'hebd8fc77f681fa3015e8efb81c8eedaa1560;
mem[149] = 144'he9afffea1947e05e143ffdb50637e026f857;
mem[150] = 144'heed4f6ce0f72e58f1cf7e765f9940988ea63;
mem[151] = 144'h0d98e715e3aa1696e87506d81010177f12af;
mem[152] = 144'h1d5aeb22119809c6f695e1eb1d9a1e161cc0;
mem[153] = 144'h0b8cef08e95b1608e2b3f897e6e4fc37131d;
mem[154] = 144'h0f240ddf072418f2ec84fd4ceaeeeb9ff32d;
mem[155] = 144'hf009e1d9faffe4cfef81fdba13c91e1309f3;
mem[156] = 144'hffb7eb15e71eeb58ffc30ea801dd161be937;
mem[157] = 144'he9a4f6011405e1781d2dfffe037419eae8f4;
mem[158] = 144'hff3d1d68ee19f732e36de2d0063d1eeef36d;
mem[159] = 144'he057f6c1f0abf982f5c911e1183919f2f7d0;
mem[160] = 144'hf050efbe1a241b63ebb61ff9fba5fb481ef6;
mem[161] = 144'h14e61d82e6c1147afcaef6a0ee0b0e62ea35;
mem[162] = 144'hf9b701811b7d0bbb02f203f8184a0d08e8df;
mem[163] = 144'h0c40e73305c4f52ce4600f27e15503ebe7cd;
mem[164] = 144'h0e6be718117b1fdaf00e1ccfe72d103c0166;
mem[165] = 144'hebcdec56f24dfaec0e9406fefe1a116df6e8;
mem[166] = 144'hf382ed30059019a01a95194e110214ab07e3;
mem[167] = 144'hedc41248f4070b1a14c702bf0be806671725;
mem[168] = 144'hef37088afbe4f99be87b19b3005be865fe9a;
mem[169] = 144'h0058f88df7700af9e6d3092e19e41b1a08b9;
mem[170] = 144'h1ae5ff75ea201501e1560e8ceae70402025d;
mem[171] = 144'h13ffeebb09390f711796f5810c32f989e3a9;
mem[172] = 144'he554e87ae6ba109b1d820ba8e5121ddc1a83;
mem[173] = 144'h0f4a0fdd19fc0d4501dde1311fc41dd30c12;
mem[174] = 144'hef4ee21eed3817a71c27fa81f360f68bebc4;
mem[175] = 144'h1ad5e8c1f4fdfb8afbe8ecc301061c29058d;
mem[176] = 144'hfeb9f331085ee8d4117dfeb1e20e1f2c1830;
mem[177] = 144'hf3fa0e43133ef89df1c3ea090e4eec21ff97;
mem[178] = 144'h06eaf4351482eafeeec20a7b01770c65f4f2;
mem[179] = 144'hf165f0530abc106fecc5155f0ea3ed4ae9f8;
mem[180] = 144'he279175ef47e07ecf2a8e70c17ad0d92e764;
mem[181] = 144'h1b961d14f31e193a116c1d72fa830996f2ed;
mem[182] = 144'hffe3f9cd1d39ef40ebc11651fdb016af0344;
mem[183] = 144'h072f0758ee9cf13a16c10625ffd8fb8be6c8;
mem[184] = 144'h1476145ae492003bfdaa0effe9fc1e040619;
mem[185] = 144'hf324f1ffe1071b661fc103e5f107f042f04c;
mem[186] = 144'h19c902c1128b17b203f80b0f12dce7c0f040;
mem[187] = 144'he8bb0dfce4270e4613c2e8ba168d195af3b7;
mem[188] = 144'h080ffe51fb49022c1e9d0470e0cff0e21bb5;
mem[189] = 144'hef5cef44163debecffcaf340119f036fe537;
mem[190] = 144'h05d3ff7d1d7af030ec53019e1ad2e43c1ba2;
mem[191] = 144'hf5c30e040f9d125717c8fd63183b09a70d61;
mem[192] = 144'h0178fef4f6da0f8306d8f8091f0ce8f7ed7e;
mem[193] = 144'h0dab1b4a1e6e03220df103671c20fa42e915;
mem[194] = 144'h114916b6e28def340bf4e7fe13bae04af62c;
mem[195] = 144'h103de9f6fcd11362e0c51586f981e78dfa2f;
mem[196] = 144'heb37e247036cf69a03e71d4fe702fa05e8ea;
mem[197] = 144'h122110cf0426e9fbf547f20200cff972e57b;
mem[198] = 144'h15fbf71ef99713cb0ac9e7c81876f1bf165d;
mem[199] = 144'hfe68f691177419c31129f298fc2df60beb21;
mem[200] = 144'h1074fcbe0a871b69e612e621fa8e1324066e;
mem[201] = 144'hf320fe80ef9bfc95153aec6fe4eae9d9e019;
mem[202] = 144'h0cd7f270e9561ca3e3711f96f13004d4f031;
mem[203] = 144'h18211b28fae511451b04004e1f73e382f6ab;
mem[204] = 144'hf43a0ab10af806adee1214a1e813e12317c0;
mem[205] = 144'hff0fe228138be765fc5e1b64e59e1b251f5f;
mem[206] = 144'h1f0aee1f1035f25cf76e0879ef7400d7e0d3;
mem[207] = 144'h1f9feeb9e9851a5be2411c32e89909a10c29;
mem[208] = 144'h093be322e3fa0aff1a4dfee7fffcfc07e84a;
mem[209] = 144'he461f168ef3109f2e5fdecfaee46f2500151;
mem[210] = 144'h1c34e08d1dd1fbc6e31e0b19fc98028b1b64;
mem[211] = 144'h0a1f140912ad13631ddae21a0bf9111f0c63;
mem[212] = 144'h1650ee4af854ebb2081bf61b197eef8cf9e4;
mem[213] = 144'hea32070010d9f3dc05481b62ea24ffcd090c;
mem[214] = 144'h14b5125900df0756e60de9c6f192e74ef9b0;
mem[215] = 144'hf5a407c317bff0ef18b6fe321afee31ee0ec;
mem[216] = 144'hf62413a0fb97fb510d7a0575fa2b1e73f958;
mem[217] = 144'h1b511c711634ec0f16e60765f368e1a61659;
mem[218] = 144'h0ed2ea7f0792f1f3f5621df1e4b40bd91012;
mem[219] = 144'hf3990431fc4c1487ef01e37e091bf3c2e1da;
mem[220] = 144'he5e6eed4fdf7ea2317b1fbfd07c3e5c0f335;
mem[221] = 144'heb65e800e7f0e2781a33ef1f031be866026c;
mem[222] = 144'h0627f160fdcdfaa400ebf19f177e153aea76;
mem[223] = 144'hee6de2ad0d811e351fd517980d0412c41d12;
mem[224] = 144'h0430169bfe011b3d06e0e7a1fb010d8818c8;
mem[225] = 144'he105fe6f0bdf127be3aef0d5146b111bf86d;
mem[226] = 144'he86aecf718d4e19b04a50b8af62efa6e18da;
mem[227] = 144'hf228084cfd2c181b15431a61e4adfd4411f8;
mem[228] = 144'h151de8d41003f48afcc8185908a701e0ea32;
mem[229] = 144'h1bf3f8b91a031d7f138ef054ef8307341bb9;
mem[230] = 144'he3a702e712c6f1df1efd10260dab06ffe375;
mem[231] = 144'h0facfe5e172e16a20ca5070ef50af464f248;
mem[232] = 144'hfebee1d61b69fac7f784f802e8761aa4e570;
mem[233] = 144'h1e49f58a19d9fa2cef21f4ae0ab1ef110b30;
mem[234] = 144'h0e1d0a07f4b0e316fd58fd451560e89df095;
mem[235] = 144'h080615aee7e51905fb1b14f61d8816cef94b;
mem[236] = 144'h1ad0ec6f0b131071ee5e1970e38ff88a1f6b;
mem[237] = 144'h118a1462f9bb05c9e7bbf0931ac9eb49e3b5;
mem[238] = 144'hf95514aff3b412ed17c106bce8f10da4e7ab;
mem[239] = 144'hf3191330e4e802bcfa211c2eefd00c00e3dc;
mem[240] = 144'h0116fcacfc50ed66fb4f0c11eeece1c800d3;
mem[241] = 144'h11531ce5ef14f2c30edfe02214b21cfef3d4;
mem[242] = 144'hf05e185c08e2f1321f9a1b87107508331290;
mem[243] = 144'h02480a33193fe599fc80e61310840e7408ba;
mem[244] = 144'hed0ef35d1f0bf05c1753f1aa067712b61c72;
mem[245] = 144'he41d1a53f76e1df2ea6411ebec7fe88302d7;
mem[246] = 144'he9320d6cf94e09a80f99eb50e887e9ff1fe2;
mem[247] = 144'h0adc080fef08fad309ae108e0288f36ae079;
mem[248] = 144'h1dbae23e0fc6001010d5119df37001ddf0bd;
mem[249] = 144'h1eb2f9ddf507e7061f8b17e408601386e150;
mem[250] = 144'h0a90006b0c7eea2d1803e4e2e8050153e0c0;
mem[251] = 144'h142b1b5ef95de38c1b360137fb2b16ece974;
mem[252] = 144'he8c60c10f62d18effe3bf409ef03e136f2b2;
mem[253] = 144'hf048e8a40fd91d5505560671faa211f2105c;
mem[254] = 144'h0976e62714fd0106e22714c60ff6ee05eb79;
mem[255] = 144'h150614cc16a81b4613f104a4eb990d1efd7a;
mem[256] = 144'h01b1e1d6e6ae01d7f84c0fd9e41d0feb0a25;
mem[257] = 144'h0b1d0270f02be766ef3614320fd3040aff12;
mem[258] = 144'hf835edf4e0b31ebaf73b1508f70e02c8e4c2;
mem[259] = 144'he3db0a81e4a50abf1f641675e33fe6d5053c;
mem[260] = 144'hff34f045fc9e1c3b1d0e0dbafdfb1161e84f;
mem[261] = 144'hf8350215f38016b005f5f39d0cc0f2030ac5;
mem[262] = 144'hf0700199ea4818bceda7062bf5f8e367e2c5;
mem[263] = 144'h03980901f6fbe570fbdcf65f0412114b10c4;
mem[264] = 144'he53cf87ff70817d6fe5a150c0b211e1af0f5;
mem[265] = 144'h0991f88ae5afe8c6f8ab1063e514e393f56b;
mem[266] = 144'hf4af1d0c0722e7e40c0d186c15010631fd4e;
mem[267] = 144'hf919f00f04c8e1d1e2a9ecbb0fb50556ea3b;
mem[268] = 144'h1fb6053e12871604174d0e0603140fbef09c;
mem[269] = 144'hf9b80d8811dee79df2bdf56fe0e7e248e21d;
mem[270] = 144'h1d30e29efea6f998002713d716811de21275;
mem[271] = 144'h1e08fd9e05bff9c41cbd18e5f0dafdc7e33c;
mem[272] = 144'hf647e73ff332ecf51c61f8e91bb4fbb90533;
mem[273] = 144'he7e202b1029ded10efa7e73f13dcf1281f0b;
mem[274] = 144'h1f8df4371e8af3ff03b2eb5b0370ede7fadd;
mem[275] = 144'h0b59030608aa002712d5016b091bfc1a1e5c;
mem[276] = 144'h02450ecce4c719251442e32f00e4f7deee94;
mem[277] = 144'h0c5b1066069f190f1c53f03502ac152a1a75;
mem[278] = 144'h18ee055f0472f84b06f2fd7b0172f7c3e810;
mem[279] = 144'h0e5718a900181bcdff7d1bf2f6071dd31850;
mem[280] = 144'h0af5f387f8181b9304011684e67ff091003f;
mem[281] = 144'he95ff5760719e7410a2d1033f7c018cc1107;
mem[282] = 144'h00c2085df6f10c28eeb6ecd005b4e933ee3c;
mem[283] = 144'h0c8ee2170423e574fd7f08f91f18ef3a19d1;
mem[284] = 144'h15bc115eeed6f35c1983ee77000af86400ab;
mem[285] = 144'hecf909c8e2eef0d410eafdda1b88e2181ba2;
mem[286] = 144'he7aeec511a4c038aefc508390d9c149ee3f3;
mem[287] = 144'hfeb703600dbfe89fe25d0ed11cff0b22ed87;
mem[288] = 144'h18ce18150180e45a1fa10e9110a9142318f4;
mem[289] = 144'h114bf9bdee381fca0d23ea841bd51f0fe46b;
mem[290] = 144'hf5d1f603f8ad04971b591cc018e10356f964;
mem[291] = 144'h1b10f24d13c0f57aff45e10c000c03ac01e6;
mem[292] = 144'hec8308d0e66e1f3c0e16e6dd02defbe7e1b6;
mem[293] = 144'he1b5fa0eff3ff5b0fbd8e95ae6a9176f04af;
mem[294] = 144'hefe8ee1a06381797f57811f2f52c1be0fd52;
mem[295] = 144'h1bc6e4b7030f14b5fe3be9121dcde65812e8;
mem[296] = 144'hf94cf46de9d1fd3ff1ecfdc91a200072ed9d;
mem[297] = 144'hec4e054bed9112f4171b028b1aedf7e50106;
mem[298] = 144'hfbd9188ae9ffe101ff3f1d9cffe71aa716d3;
mem[299] = 144'h0a7e0e30f3660f58fb5ce0deea1703ec0fd3;
mem[300] = 144'h0c0af8a1f541f4fa09f4eab009efffe6f811;
mem[301] = 144'hefddf5bc1779ff3bdff701dafe32e44d1a0b;
mem[302] = 144'h19c40b101aa1e21f1178f99ae783f19df4d9;
mem[303] = 144'h189cf255e7a8e234f9be0e9c1d22e2060ba8;
mem[304] = 144'h10091bfbef3d145eecab16990b5412fc1603;
mem[305] = 144'he656ebabf91d07a8eef304dae53e019debe4;
mem[306] = 144'h19951342f9930727f0b3ecd215dd170ffa42;
mem[307] = 144'hfddee63bf48d05abe85ce84501ed16c3f277;
mem[308] = 144'h1a821e6af5851cf5e7d016fa0c2d1f261903;
mem[309] = 144'h18b8f4bcef2717fff0d31f95f710e3601a7d;
mem[310] = 144'hf7d60bb014891a6e08b5116c0c4ced031359;
mem[311] = 144'hf0960967feba1bb00552f686ffd61c85f0f8;
mem[312] = 144'hf8dcee7e0a820986e9c3fbf7181bfef4f6a8;
mem[313] = 144'h1c3dfffbfda31afbf9e1021713f4ec1fe128;
mem[314] = 144'he41715eaf071135509fc1b6ce67907a7091b;
mem[315] = 144'h06fce2d2ef4c14901e73ff02e8701d7b00d2;
mem[316] = 144'h1b6de000e8dfe9c21855eac81e84192e1764;
mem[317] = 144'he22d1120e935efac1e57e9261cb4054bf696;
mem[318] = 144'h043b07571d22fcc90987fc8df5cd02f0ef75;
mem[319] = 144'hebb802d0099ff445e697f8ed1d981485e39f;
mem[320] = 144'h0ee7e7f0e43cfce11f7b1989137efd20efe5;
mem[321] = 144'hfca2e88affb20f13068201c31ab2022f17d2;
mem[322] = 144'hef29048600a619af1540ede4ef8ae04b1e50;
mem[323] = 144'hf7981532024df684ed9405f30f3e1a5cec8d;
mem[324] = 144'hf219f530f2b417f3e54ffb270409195b0e23;
mem[325] = 144'h1aa60fcb17caf1381b82e37d17fcfed81b40;
mem[326] = 144'hf3b7f5601f941a4700c303a416bffb7df9d7;
mem[327] = 144'hec020796158108b80df70336183d181d07e4;
mem[328] = 144'h1f2018a4eb711150edee07cbe722ffbaec77;
mem[329] = 144'hf004023413eafc280421e514f0a2f39ff479;
mem[330] = 144'h0fecf689fdfaefe7ed2ff8f2e6a20fbbe8cf;
mem[331] = 144'hfc24036cfb90eb950d46f5ff11c106031ccb;
mem[332] = 144'h048ae6d40e20e59d0db9023be1b7fc85e49b;
mem[333] = 144'he2860e1ff6d4ed72fdf11149e9bb0ee4f2bb;
mem[334] = 144'hefa9006318ba0e17e82df19c0a0706cd1351;
mem[335] = 144'h179217f81451fe8e1304154af52ffe73f1ba;
mem[336] = 144'hfb9b04d91d8e13fe1c97f053ec34faa9f756;
mem[337] = 144'h0bd6ef5ee07517b1e5e211411b3efc031f44;
mem[338] = 144'hee14140c034ef959eb35e08bfbe1e801ef3a;
mem[339] = 144'h1ab6f429176eed3b15310e32f192f67cedc9;
mem[340] = 144'h1cdefaed1ab0ea6215b40400ed0c0f12ed0f;
mem[341] = 144'hfc0713850201128eeb6a0fcce75b1521f26a;
mem[342] = 144'hfb3e0c21f5ed185a125d17a91a770038104e;
mem[343] = 144'hf14dfb8becae1f2301831cbaff7503f2e35f;
mem[344] = 144'h012dff30187cf65d0ac91a500bfaf4a3009a;
mem[345] = 144'hee29ec0fe17ff69f00c0f619f940e687fd5b;
mem[346] = 144'he4f11075eede1a3d1ea2e1f3ff0d11be128f;
mem[347] = 144'h1ec5e3a3024d15511a8fec290e241c7b0e4c;
mem[348] = 144'hf270e5ee10d0e71def550f92e3aff4830feb;
mem[349] = 144'he655e537148cff72e5b10c16e60d035d1ab5;
mem[350] = 144'hfa250f07e9cf193ef1ce187ae837ee4ee398;
mem[351] = 144'hf010fd8ee472f10ce153fa2ae33801f4f966;
mem[352] = 144'h16ecf2930c4bfc37f10d03620bdd1b310082;
mem[353] = 144'h12a40b3c0f2a0a2a19b908c50e25f49fff10;
mem[354] = 144'h1f6ee5841d5f0c56184ff33e1509119be6f3;
mem[355] = 144'he0be06520231f0c7f4b9e25fef3cf7d5fc03;
mem[356] = 144'h0bb9febf004ee963f66f0ee5f803ee20f5cc;
mem[357] = 144'heeddf9310ecb03c91f84f39a18231b1e1c40;
mem[358] = 144'he82f1e68e00aedd2003bee6117b5ecd1f5bf;
mem[359] = 144'he983ed3ee8ba0846f3500b920dd5e9540f2d;
mem[360] = 144'h0a14e29ae0c70890f0591160fd060c740c15;
mem[361] = 144'h140d1b231f601018f0c60c600b8eedc3037d;
mem[362] = 144'hea60fb28e392f11f1af509e817bdfcdc0472;
mem[363] = 144'h09231981055ee27106c20232ee190458ea84;
mem[364] = 144'h06ea10a40133153e1ea5eb7d1e28e48de314;
mem[365] = 144'hfa411322eaa2e33310361804edd1fdd1e56d;
mem[366] = 144'he298098ef82ffef419f2f077f4b106831a4b;
mem[367] = 144'hfd9d170e054102c40ab0e82e1282038714bd;
mem[368] = 144'he2bce5810abaf549e6b90a49ef9c031818c7;
mem[369] = 144'hf10b03870717e1390084f2d8e90800190f8b;
mem[370] = 144'h1cdfec4c16bfed16f1e6f191e9c6e14e1334;
mem[371] = 144'h1b79fe0012cbe6500f48eb4610a3e68b0449;
mem[372] = 144'h078c1a3b0512099619f61d7f0860e46d062a;
mem[373] = 144'h073811a3f9c9e3fa0e150bda0db013721428;
mem[374] = 144'h11b80d2be409e0e7ea8513cb1151082af603;
mem[375] = 144'hea8608f3e224fb76f9bcee1df8660e42f59b;
mem[376] = 144'he7d00d86e3b0eac5e68817cf1621f1bafcf8;
mem[377] = 144'hfc3b10b9fb78fed014f7f1c6e073f524007f;
mem[378] = 144'h141018fe01881cf5e76e12b7e603e3e1e7d2;
mem[379] = 144'he02b01790813fd08105eeda5ee65eba9ebdc;
mem[380] = 144'hfd7a129209490a13f0ef0f2ef56c1af9ef34;
mem[381] = 144'he69ce34813c00fd803261493fa5cf5f51446;
mem[382] = 144'he33810181e91f72e1b72f4d509ff15d2031f;
mem[383] = 144'h1430e3c6ef8efceefee11b10e687f4480305;
mem[384] = 144'h019e1ddde12d1d0ff90c0c73f9c6e5eee32e;
mem[385] = 144'he372f759f58a1120080110d9f51cea551092;
mem[386] = 144'h08d70846fe83e407166605931098e92ae2cc;
mem[387] = 144'h0c620a210585e99bea3eeeeb1d730a181a99;
mem[388] = 144'h031e049ee34f129104fce3c900f8e5ab0733;
mem[389] = 144'h1bf3005a0dcc06fe01ed0922eb091f2d0196;
mem[390] = 144'hed580656fdd2e5e40069e9620ffae12f072d;
mem[391] = 144'h131ae34e122bf1c2f58e0a1e192ae5ba0b9e;
mem[392] = 144'h07fd08c31144f1730af0ea9fecddfd991dd3;
mem[393] = 144'h10b81861fd7f0448fccee986fca608a30a96;
mem[394] = 144'h160fee4a1ad0f6881c171d530c62f4fc0537;
mem[395] = 144'he5750e2d0db2f7c0f672e19904c60b45ecf7;
mem[396] = 144'heed5fe6f1a870e55e42a0a3402a011dd1daa;
mem[397] = 144'hff1ffa4508a6014d189ffb9ae527ffadfa38;
mem[398] = 144'h0f540e171f670ede0198e7f0fd65fd53e19b;
mem[399] = 144'h0caf0c93f82d12ee05c0ff3be77d06c1f2e8;
mem[400] = 144'hfd220fa005da1e2b0adc1d91e8030e94f3b5;
mem[401] = 144'h12d6f89ff92d0e7a0b09ee0e0980e1560937;
mem[402] = 144'h003be411182c07cd139ff95e180af46c1d54;
mem[403] = 144'h148df0b41866f48a0ecf0dbaeaa0ee01f438;
mem[404] = 144'h11cafb31f113e4a1e345e7a7e83ef0cce435;
mem[405] = 144'h0830f86a0cd31089f199e7b1194f03d613d6;
mem[406] = 144'h129aeaf61f2f0df214a3052d0cca14371c33;
mem[407] = 144'hee150dda12cf14f5f1090b980f2100fdf496;
mem[408] = 144'he6a91ce5e2f6edf6ebfa192f0a560bb410be;
mem[409] = 144'he9c1fdf20ae1ebf2f88e06e1e5b206ad03f0;
mem[410] = 144'heeb704affd2612c1fa3a0384e85ae162f202;
mem[411] = 144'hed90e8c1ffe0fb430df9f09be209fe50e27d;
mem[412] = 144'h1502f6190d6708c4f711146d1905eca41a73;
mem[413] = 144'hf7b7156ee8dbfa05f0bae88de779f199ef8f;
mem[414] = 144'h0b3fe433eeda079de1b0e12c036f035815ce;
mem[415] = 144'hfbe005c719df0dc2ee2ffa521958024b07ea;
mem[416] = 144'h15c1e876f977fae6f848facd0536f5be00d2;
mem[417] = 144'hf019039b048003e8f1f9184de61005770282;
mem[418] = 144'hf6eb0f8df8f40c09ec1bebee002319e7134e;
mem[419] = 144'h16e5f236fc5d060ae3701151f83b1774f1fc;
mem[420] = 144'heeedfd15121befa6edcde85f151ce9b1eb4d;
mem[421] = 144'he382f880f3081d44e808fbe1e4f2e4150c95;
mem[422] = 144'h169415f4e288f3bdfb72f890064ff59eeb57;
mem[423] = 144'he4470c3109d01b7cfc16e46d178de12cedae;
mem[424] = 144'he2610a5b1816fa84f757fa440266ece0e0db;
mem[425] = 144'he5e20568f3f0f9fd1272030e0166f4340da0;
mem[426] = 144'he84be8d5fe0ae608ef2a09e60d1b04091b7f;
mem[427] = 144'h1a65f0c0f1b8e60aebc116f7ff64e7871bc2;
mem[428] = 144'hf1eb0f70f0ddfd93f4e81c5314d00d1107f2;
mem[429] = 144'heff01e7b041f05541ad80837eb6104d7e513;
mem[430] = 144'h0cac1c08ede01b4bed7feac9eec60ba1fcd0;
mem[431] = 144'he350153e0210ec85153ce682f5ee086ee003;
mem[432] = 144'h18bcf27b18181f9810a610c6eb4114b40a3b;
mem[433] = 144'hee64f4d30b0f15f7f6bbe9d608e9f186f87d;
mem[434] = 144'h112e069de325f2ff1ea1f924047f074c1d7a;
mem[435] = 144'he7140c3ae5f6e9d70db805b8e632f92d079c;
mem[436] = 144'he7761ce1026fe0afe963136015b9f74eeb1a;
mem[437] = 144'h1f3f1873e528e46fe87cf1e10ccde56f17f8;
mem[438] = 144'he053ff5cf776eda3ea1809960b78eb56e786;
mem[439] = 144'hecb6e3f10c4a1d18e69ae6c6efc3e7d30a69;
mem[440] = 144'h035cf2041134f22102c808e9ff38027719b5;
mem[441] = 144'heb3cfe0ff96af7c2f6f0e646f918e4f41e21;
mem[442] = 144'he559e66bf8f10abbe1b0ee3ffd79f3b1f7c1;
mem[443] = 144'h0d5df03ef740ff861d13f0efeeb91a49e604;
mem[444] = 144'h17c9e751e5faecbcf472e6bff2efedad1ec6;
mem[445] = 144'hef870a9106191759f12119731ed3e9dae65d;
mem[446] = 144'h0752ee710819f732fda5ed6bf52cf36b0170;
mem[447] = 144'hf56112961bfc0c9cfed0f0b3fc34f0bde134;
mem[448] = 144'h19e10922fe46f86afbe9e5b0f80bf97f0d53;
mem[449] = 144'hf91ee9b806e40d64e8c00af40765069d07a0;
mem[450] = 144'h12331319f3ad0494f03de9e5167de1041102;
mem[451] = 144'h0d1f1e4d1b7de402e7ca17de1bd0fd0cee1c;
mem[452] = 144'hf69f054f1c25eee2faa5ea40f4b40b9616d0;
mem[453] = 144'hf2ba0eb90798ede90fc7e81e0a791e240454;
mem[454] = 144'h14b0f09deae2e77f0b2e0301f32ef175fd5c;
mem[455] = 144'h1aab07ffe2b2eaafe94100111ba0e64ae013;
mem[456] = 144'heaa311d8e640fce8e668e775f35bf89d00e4;
mem[457] = 144'hed520f4812afe652e4300c1d1f3400621aa0;
mem[458] = 144'hecf8fc3a1f01f141070c000f00c4fc81e1fd;
mem[459] = 144'hf64e12aff39afcc50de50d66e68612731d97;
mem[460] = 144'he6b2f73a0471e622f0260eda077e0c751e09;
mem[461] = 144'h15c0feea1e21e1fe1eb9114607c113e2e624;
mem[462] = 144'hfb930e10e9f715ed1482153018521bda0eb1;
mem[463] = 144'he836eed210deea8e0367f49ce10d1f6cf7ee;
mem[464] = 144'hfddc0637f734176d04d70549023a199b08a3;
mem[465] = 144'he0f41e45fe901e9702b2f14ff3320a071493;
mem[466] = 144'he1daea48f47ff43d11d415441f06f3f206ea;
mem[467] = 144'h034ff216facae0801efbfd121363eba3eb03;
mem[468] = 144'he660f90d0268f050182a01a2ea23e6890517;
mem[469] = 144'hef4810e3fddc0fd8f5d202790bfbfca40b64;
mem[470] = 144'hf233ed0f1777f740f18ef895029c0b621e7d;
mem[471] = 144'hf2ff12031bd1eb8d16d80675e1a3e91e101c;
mem[472] = 144'h1264e49efc840fda02c116151ca612e30823;
mem[473] = 144'h01aef1e10cfc1b77ef6af3df0a1a030ff888;
mem[474] = 144'hf4190b6fe3cc13951aa7080c186d00bc1a3a;
mem[475] = 144'hf05d191300b90debf99b0f6a1a6102aae00f;
mem[476] = 144'he961152903c3f4bce2e9070819a8e0bde5e5;
mem[477] = 144'he0b60f7ffbc112b9e540190ef5a01a4df899;
mem[478] = 144'hf51017aff77a0133f53e01a812071791e5c0;
mem[479] = 144'he2ed0a2a0ad81ff8f6de1e2d1233e7ea158f;
mem[480] = 144'h0f7f0b400f4dea09f3f8e614ff80fefaff17;
mem[481] = 144'hecbc014c155e075ceeece4e9e2e6ed5013a4;
mem[482] = 144'he3580f2efd8213cf13e1e99312a2ec591f5a;
mem[483] = 144'h015016a601b4118d05f41ef80ebbe450e10b;
mem[484] = 144'hf86003b8fa6e1a61e5f30d5a16dc18c6eceb;
mem[485] = 144'hf91b001a1d650af3f809f5401e89198ce22c;
mem[486] = 144'he7001ab508d8f55ff804e94e1b55fca412c9;
mem[487] = 144'h0115fcbf06501cc3045ce4db123af50e0f33;
mem[488] = 144'he898f2970528eea201221a5ee508ea9e0e17;
mem[489] = 144'heffde83c0fbc103104471b46053e0fcaf2a0;
mem[490] = 144'he183fa68126518b109bbf659e25718efeab8;
mem[491] = 144'h1258fe4beccdfb1b1074f44804860fc306ea;
mem[492] = 144'h0dc31dc306e6f0a4e2aff47b195415cbe1e2;
mem[493] = 144'h1ed9f39109c7f0e4e6ce1eda1648e5dde28e;
mem[494] = 144'h1387ecf8046217d21378eab2faa206e2e273;
mem[495] = 144'h0ca20c751b45f3d9f3861dc20a1ee7910385;
mem[496] = 144'hec2714261f52f665027a0cd31c3ef1aeeadd;
mem[497] = 144'hf80710c1fa5513dd01d50f66ef9c1d6c0a4a;
mem[498] = 144'hf4b31073ff3df764ffde0b7ef671f1a10401;
mem[499] = 144'hf41419af0c380ba7f140f0a312dc1236010c;
mem[500] = 144'h1e971f241db4f7861b831f63f451fde70b3a;
mem[501] = 144'hf091fa26f56e0449fa2fe406e3a31a6f109c;
mem[502] = 144'hfacb118a18c606f6f965ee740d27196cea0d;
mem[503] = 144'h1ee4ea1be8ec0874e67007c1e9e01349037e;
mem[504] = 144'h120ef53106d7e43a075fe9f2f5a30aa0e193;
mem[505] = 144'h1e8e185304c0e5c6e65511ee10d01be2f19e;
mem[506] = 144'h112ef4bef870e175081e055016c6e71afae6;
mem[507] = 144'hf4e20655e5870c05e8f10eade7161b001dbf;
mem[508] = 144'he3adfa76ea6aed24ef2f124de5151453e318;
mem[509] = 144'he6430fb5ee4c03d709f3eeba17a5fe2cee33;
mem[510] = 144'h17d7f453ec61feaced860c2ef68fe481f617;
mem[511] = 144'h114ae649f44afe0bee45e0fae0e3fe86e0aa;
mem[512] = 144'he98816c2ff7afa7a14b015f4f45e0a51e902;
mem[513] = 144'h064fe750f8e50c351df0e566e368fcd5ec88;
mem[514] = 144'h132518620d380cb71aa10ff40019e1a2ffab;
mem[515] = 144'hea53159de37de7b6fba00c2b04b3134fe027;
mem[516] = 144'h074e12270658e26f1be50711f142023be65e;
mem[517] = 144'hee1017660c20e9781585e63c074b1d67eb63;
mem[518] = 144'hea21133d10f3e0b0e8d0f3c0113df22b1290;
mem[519] = 144'h01351b19111502f00863f221e47c1e351fb4;
mem[520] = 144'hfa83ecf3ed37e46eea49e99100b2f43c0adb;
mem[521] = 144'he2b2ef6707bcf61003cb023a12d0e01b11bf;
mem[522] = 144'hf14e1e5606ca0aaaee1ce9daf8440cfdf673;
mem[523] = 144'h0eb9fbd0125101dde628fc910a610a6b0c17;
mem[524] = 144'he12002061fa9fba40f11e4180774154e0af9;
mem[525] = 144'h1e8cf32006cf126217c31e6416030da816af;
mem[526] = 144'h1276f309138cf6d41125ed7a19e007f51fdc;
mem[527] = 144'h0701ed2f1800fb8c0606e0e7fc1d1bef1195;
mem[528] = 144'h0ea7ea57e7c50df1e8841399e45f07951c59;
mem[529] = 144'h0ff809d31c181e94e083fd95eeeae5a4fe07;
mem[530] = 144'h0855fb76f781088ae676e0f3f0541528f033;
mem[531] = 144'hf4761025f5c90e081b8d0631f726fda80395;
mem[532] = 144'h04dce5a51c3e09a7f0fcf2a91714e531e043;
mem[533] = 144'hf7f8f084fe0f1e0c07a8fa61ff0711f903f2;
mem[534] = 144'he38fe83cff0fe5aa1de8e6f604fc03b70de6;
mem[535] = 144'h04721ced076b0965fee4e29e16fef7dcf86f;
mem[536] = 144'hf455059de9d3ef63f16c0e842010f5b010bc;
mem[537] = 144'h124814e9ecc5f0e9e8b9fa1f1a89eabcf8d2;
mem[538] = 144'hf2f50b16032f0df40367e518e872eb18009c;
mem[539] = 144'h0921fe7affa3e344ec701373ee94ffa61c34;
mem[540] = 144'hf505e260f64d12460f0af4c31bd410cb14f4;
mem[541] = 144'h0425f685eaf4e9e1ef25e9f4f1e31ca01f05;
mem[542] = 144'h1b3be28df04fe3cae726074f0f90e7c21aa7;
mem[543] = 144'hf921f967f162f5540c7900f1e8aae88a1812;
mem[544] = 144'h154e0e63008a040e0a1cf960195a0a54e753;
mem[545] = 144'hea6905be1930e586fd5605a80b5b1bedeb1a;
mem[546] = 144'h1ee6ec001c411dbce8b1e91b00a210eaec8b;
mem[547] = 144'h0af3f09612bdea5c0081f1e1ea53168e0391;
mem[548] = 144'hfcc8f83910b4143fe24903421347e8de03f3;
mem[549] = 144'heafee0ebf0371f81eadf0ea7f3771c74020f;
mem[550] = 144'h10fdf556e46203851d81f65e1d9ef310f38f;
mem[551] = 144'hee42f8b704f41f5f16a3fbc102991a4d1680;
mem[552] = 144'hf91403e8006113e512c102b0ea46ffc1e81b;
mem[553] = 144'h0ddbfb9f199efeb30fde136ff3b91aaa1687;
mem[554] = 144'hf1f6f023024ffb99fe0e05930a97f1c3e1d5;
mem[555] = 144'h01aaea1d03c7fddefd280bb01ffde98fffcc;
mem[556] = 144'h0b81e050fc35f78c13f3e1930d3a1311f4ce;
mem[557] = 144'h1c19f1ba1d3e13fd03a21a5e0634ea47fb44;
mem[558] = 144'h1595163e1a90e7bafec2057c1775fc84e42b;
mem[559] = 144'hf7e218d5fceaf2010e56f280eb25e4971068;
mem[560] = 144'h1e9f1163eb10f668107ff67c08450ac915eb;
mem[561] = 144'hf8a4069803371f7c0f26faedf3f71dfdff9b;
mem[562] = 144'hea21f365f12aecda16efe1f7e5080e28ff89;
mem[563] = 144'h01891c9ee06be7b1e41af1df18bb080be4b8;
mem[564] = 144'hfc881140e718e55cfddb029bf0cce20ef6d0;
mem[565] = 144'h112be63ffe8cf36be5c61610e9580b76f377;
mem[566] = 144'h1718f5b401251df6e0e6f7e6e1f71c7ce930;
mem[567] = 144'hf7bb17b90073140b1af8ea9a013b09051d35;
mem[568] = 144'h19a0e051fef61b9bfbebe834eaf707440bca;
mem[569] = 144'h0f51fa65e645ff990762eaceeab0e55a1684;
mem[570] = 144'h03870ac3f3ddebb60574f736f18a0dedee29;
mem[571] = 144'hf14df2daf9341d73ecc4ff9606c7ef5d06a4;
mem[572] = 144'h14f60d580be8ec120adafe2dfd0af913fdef;
mem[573] = 144'he9cbefef1dff0bad1fb6f378ff94e8d11ea5;
mem[574] = 144'hfc6fe4cf18f6144d02d8e31212200d5eece0;
mem[575] = 144'he50a1124031c08cdf4eff18dfe9a1dbdf154;
mem[576] = 144'hf10f1884e5aff2a201b40bf31f08ee580252;
mem[577] = 144'he30c17050565ec3818eae941e2261011ec96;
mem[578] = 144'h0778f4870fb50649e13213c2e39414a50d7f;
mem[579] = 144'h06e61637e3780b980a2f0bc319baeb8df967;
mem[580] = 144'hfa14ecc3f240e0bc056619a21987f180fba6;
mem[581] = 144'h051a134e0729e371efabfa251d0a0d7b0cce;
mem[582] = 144'h12aaee70f9ff10ed009af26a01d210671f8c;
mem[583] = 144'h005c0f4d15351a75f4d4ed7ae8ebe57cebca;
mem[584] = 144'h0a770c39e7dff623e891155eea07f2e70d5c;
mem[585] = 144'hfaa418cff2e81aee0f780f5a1691f693eeee;
mem[586] = 144'hff0eed0418ff10ed01bbeda2faa0ea6d0bff;
mem[587] = 144'hfdbf060f1f0e0b0312f5effc01ce1e4b100a;
mem[588] = 144'hec11eb320b490dd91bbe0ae8143d187ee63e;
mem[589] = 144'h018a11b6ec61fee6efb118b70f83fa5b06e3;
mem[590] = 144'hf888f274164706f9fe77fb7007b0eaa0eb9d;
mem[591] = 144'h07fd0cdce4bdfeff0fe2e47819751d501c6e;
mem[592] = 144'hfa59180a19bfff03ebd5ee86092aeb7cffeb;
mem[593] = 144'h0f84e7cb1adb02db1905ef2e10670f400334;
mem[594] = 144'hf3d1fc681a32e5600ea4e30908b011041f3f;
mem[595] = 144'h10ac15edf18de947fcc213f11092e1f0116e;
mem[596] = 144'h1982f699ed9bf7660e83e48ae80f10aef18a;
mem[597] = 144'hf5131ef1fcbe1d8ae6170cbd1e5ae8761d2d;
mem[598] = 144'hf2fa1fc7053bf673ec711c8df0fc0523117a;
mem[599] = 144'hfd971db4f5e903d61cd50b8ce50f01a7f1c1;
mem[600] = 144'h147bf32ff334fb4ff188021ef22ee33f0e71;
mem[601] = 144'h0184f3d41971ea7eea23f218f221f1a0f283;
mem[602] = 144'h1082fc07ec60ea390fabe4cbfb9e0c820bf0;
mem[603] = 144'h204613d50d16165204511dd41a4919d0ff6c;
mem[604] = 144'h1be60a66f1f215430573ee8fe9a516f5e9f5;
mem[605] = 144'h05eeeec0e8c9e25cf1bfe5b3eef5e12b0ba8;
mem[606] = 144'hecb5e2abf3931b0be80f1698e2ea15421ca8;
mem[607] = 144'hf0f3f9faf35dfc91e3d5e4cb0bf2eb42e228;
mem[608] = 144'h1f801d47f13c171fe34aea5b1bfc09120262;
mem[609] = 144'h07540f1df82914220800ff6fe9c3f7fbf485;
mem[610] = 144'he56ff721056802d714420aa20777e7b7f569;
mem[611] = 144'hea7c11bcf6e0e3b3e96be4e0f727e84e04a4;
mem[612] = 144'hfaa5edeefa8cfa6bf5581ef616d11c14005f;
mem[613] = 144'h1949ffc9e55efb6deb45fb9717cee61a02d6;
mem[614] = 144'h1751ee911dd91ac016a01edbeca9fbe200d9;
mem[615] = 144'h1b3415421838f4030ef409efed22e837eb9c;
mem[616] = 144'h1723ffc5e8b4ff750a04133e0ecf13351547;
mem[617] = 144'hfb240fea11bd15b1ebe1ef8eec36ec7ee9ec;
mem[618] = 144'h1cdf1602ecf4f9550791fe541379ee1f0089;
mem[619] = 144'h1eb51b9bf1551428e0dafc13e9320de4e1db;
mem[620] = 144'h00250ec6e9671f01148f176cf249054b0dc3;
mem[621] = 144'hdff6092bffc7181ff232149c14f5f4d71808;
mem[622] = 144'h00971969f0ff0af4e4dffb021fd01343e98b;
mem[623] = 144'hed41e4e4e8d1ef61014c174ee5dee04beb65;
mem[624] = 144'he99bee8bf1f618f9fb1ef14119f7e0ca1f13;
mem[625] = 144'h1f8b1f8e05e71ac10a801d201b1f1dc7f593;
mem[626] = 144'h182408111a061628e76ffd35e53af8acee21;
mem[627] = 144'hffa5fe5311ffe8a3119ff7aaffc4f433f9ce;
mem[628] = 144'h0b88e036001bfaa0e41319f714c8e0fbf0d4;
mem[629] = 144'h196efb8e1e12edd0eb85ed1b0fe2e7a6f095;
mem[630] = 144'h0efef16c1d9a1c9b16501adeeb9513d9f834;
mem[631] = 144'h0e06f9b3f3d9fc6de563023af63fe3001be2;
mem[632] = 144'h19e2f9bce35c17d1ffdce50e0adaecda066d;
mem[633] = 144'heb7c14c7eb3a11131bcef0cffacef6e11ed0;
mem[634] = 144'he7b3e0840ef0185804970e120db002f3e183;
mem[635] = 144'h0b4c05aee0320fd20dd1fa120277ec0fe42d;
mem[636] = 144'h0996ee2ce25713f4084af6e00f3af3b8041e;
mem[637] = 144'h0945188efcfa00cce2bef38cfec9f5b7e772;
mem[638] = 144'he374ecbee17fe1591543ef0ee6140814e5b6;
mem[639] = 144'hfcccebd9e982f765e63b12870658f3e5f306;
mem[640] = 144'h13c1102202050228f1e8f34609141b9ef528;
mem[641] = 144'h135aea2503a4fdc21090e716f68bfa1cfe7a;
mem[642] = 144'h05c71c07e39fe299ff38135b06e3e1cef61f;
mem[643] = 144'h10ef1679ec15e0f201fe13980a270ed1017c;
mem[644] = 144'he24dec4415d6fda819111c18fd0ce41de05f;
mem[645] = 144'hfb7f0d09eccbf3f4f2d90d69f773f7a3e12a;
mem[646] = 144'he3e7f64c1fe6f5430491f0bfec0607caf10b;
mem[647] = 144'h0af200500bb2f0fff72bff24045cee550b79;
mem[648] = 144'h1c470820f8980b65f8a4ee22ea40fc011e70;
mem[649] = 144'h039000931b280273f15af788e66ef2981535;
mem[650] = 144'h12ab061cea0a195df4ceef77e80a1ff30d6d;
mem[651] = 144'h1a9518450a151477ed3af3d60339f05318cd;
mem[652] = 144'hf3bcf45217b0034818f209e3fa8104511049;
mem[653] = 144'h191e10e4e302ef34125707f915d719d0efd0;
mem[654] = 144'h0e471b44023d045e0ec209b40f881adde5fd;
mem[655] = 144'hf4d106611feeea7eeb2bf6c3f4eaeaabee7c;
mem[656] = 144'h0a5013bce52e1d98f31916e3fd84fb24f471;
mem[657] = 144'h1707fef01c8608ef08f801250f83e6ebe269;
mem[658] = 144'hf35cf25c03a2f513f63df6ee02d7e00be5d0;
mem[659] = 144'hf3411b78fa04ec1be5a01d55f27c1179f91f;
mem[660] = 144'heb66fcd111e5fdd3150e0b00e8330ab51b33;
mem[661] = 144'he496ed85e57b1bcd07dafa1508211dc41035;
mem[662] = 144'h0a9cf78200def014f428e496f2a8f70b0632;
mem[663] = 144'hea570937e051e90ffb09e16a1545ed59f602;
mem[664] = 144'h098409830f56ffbef7aa16d3e1c6f83e19f4;
mem[665] = 144'hf295f44915dae93817a3194ee082e5710666;
mem[666] = 144'he24e1bc311d1ff7504f8ec01110af145e631;
mem[667] = 144'h1e17f262fea80be3e783f713f42d0048f6fb;
mem[668] = 144'h0210f1fdf693e062105408def9c80cf5189b;
mem[669] = 144'h040f1788fa70e21ae671fddee087f11f16ad;
mem[670] = 144'hf10c199de9111517febee486f5ec1972fb5b;
mem[671] = 144'h1e8203f106d31d1c0b49e3210dc5fc7feb80;
mem[672] = 144'hec98fc7f047f1a02fcb1eccaf259e5b4eff3;
mem[673] = 144'h0b95fa3b1abaf289feebee681e40f874fbbc;
mem[674] = 144'heac2efa8e0310d661187e19f16c7e073086c;
mem[675] = 144'h15b0e18d0c6ae48919a11f99e928e982e44a;
mem[676] = 144'he6030ba3055b0315f7de0e80e5430405ffa6;
mem[677] = 144'h094ee4e702c11e4310e11ac10d77f734e081;
mem[678] = 144'he4a5029c0e35fcb7f8c1f587f82ae3c0e6e8;
mem[679] = 144'he90c1189f59211171f1718731caf0493fec5;
mem[680] = 144'hf88ce41f09fa173d17b108041b5e028ee3e3;
mem[681] = 144'hf08013fdec5e067c07b51656e2b6e7f6fa52;
mem[682] = 144'h1eb9f25ee20af661e30ae35201981e6fee2e;
mem[683] = 144'h179ffbc718ece4fbff77014bf42b0a84f7ce;
mem[684] = 144'h1c2ffa221b2ae733127ae8ab1a70f9ab0349;
mem[685] = 144'h02a3faca1c741cda15891988e7b6f4acf538;
mem[686] = 144'h07c51fcf1b57ec78e448e97de3e61797ed7a;
mem[687] = 144'h09f1f131e3c9139816a5f6020189e31dfa94;
mem[688] = 144'h0a9405d1f909f7eff287e1e11987e4241bd7;
mem[689] = 144'hec101b250971e203eab31cdb02d2fbd7e0d2;
mem[690] = 144'hf5b81ae8e9c8170ef23eedf3091ceaaef82d;
mem[691] = 144'h0b800ea81514e26c178ffb3bf3b612ed11d3;
mem[692] = 144'he803fdf50137021810fde5faeb26ef23ee26;
mem[693] = 144'h1595fd3eea51e5b8007e08b0e2ca1b48f0f7;
mem[694] = 144'he603031ee9550f5a10b6182508840fea0bbd;
mem[695] = 144'hf5861a5afd4406f011c5f45702a4fb80ffa1;
mem[696] = 144'h1bac08011d51fed309110d370f74f92d102d;
mem[697] = 144'h0623177cfdbe19a6e4dc011d04c0fe08eb1b;
mem[698] = 144'h00481501fafcf5cfe989fbd20f340dcb0229;
mem[699] = 144'he263fe58e59ded31f85ae6e610a90a37e7f9;
mem[700] = 144'h0ed9e545036de294f8b0ed4d1006ebc31c32;
mem[701] = 144'h1808f097f52ae6cb117b16e0fd8705390ecd;
mem[702] = 144'hff1116a8f502ee6a035ee0e1ef53e36d0325;
mem[703] = 144'h0078eeed1cecfd3b0e40ec4104c11eaee737;
mem[704] = 144'h1259fcf9f498ea3f0c86e747ea8111c1e1cc;
mem[705] = 144'hfc24e2c3f3461b0403b7ebbaf615ecacf4bb;
mem[706] = 144'he44b1b3ffa14000e14bb0d7bf150e9a018ca;
mem[707] = 144'hf505fdd802f4f3b4e39afbb8f63cea9510ea;
mem[708] = 144'hec11e837f324007efbfee8ac0e8f192218a5;
mem[709] = 144'h1986f88ce04d1dcd0bc6f82b03bce5cf0321;
mem[710] = 144'h010ae6d0ebf5e6380b73e077f8521ff0ed33;
mem[711] = 144'he0c20cfef287edef036b093b18e1ee01f833;
mem[712] = 144'hee17ff4f0056e32efcf9e71c066cfb920050;
mem[713] = 144'h0c12f246f2beeedc15f1e6c5f09b017be4a6;
mem[714] = 144'hea8be8bee9de11f302f6ee90f64e10c007a2;
mem[715] = 144'h125000731cdc1222f60fec92ee741b731082;
mem[716] = 144'he6fef7080fc6e4610e13e818fef202e0fd52;
mem[717] = 144'h0edfe1b503ffeec7096ce235e3a4fd65160a;
mem[718] = 144'hf6a10d82e40602a2ff7efbc206031d71fe03;
mem[719] = 144'h126c0c9901ede987e60c0b9802a101560fe0;
mem[720] = 144'h05f50cb0f3681d431d35ee59f22bf41606ed;
mem[721] = 144'hfbbeeada05c8f5ce09be0a0e13c6157704b5;
mem[722] = 144'h09ddf3e4eef31faeeb1d0328e6eb0105fb50;
mem[723] = 144'h027505d81a66010308f9f5ade8f10de70467;
mem[724] = 144'hfdca13700c2b11fd012b13e2ff2bfd8be7b4;
mem[725] = 144'h0823ef4802b70737f40af7260342e832e939;
mem[726] = 144'h0ed7ff11ef371220e830e995fdc2058018db;
mem[727] = 144'h033a07f71138fe1c087b13ea13fcff14fbba;
mem[728] = 144'h111ae0bf08b305cfe1081b1df74eea6beb91;
mem[729] = 144'hfedfe6150b8e06970e79062d0132f5c31de7;
mem[730] = 144'he38212c400731a60176ffc571fdbf5edfbc9;
mem[731] = 144'h1eb80169e5b6f70f04edfc38fa3f11f0ea5c;
mem[732] = 144'h129c148c00f0eabaf52713c6ef651b501804;
mem[733] = 144'he76018c91963f86b111111a702ea00eaf276;
mem[734] = 144'h0313fa721c26e74a1fce1687ec7cff8de582;
mem[735] = 144'he78507de1ae6f49d1c400e97f421ffaff567;
mem[736] = 144'h0da010aef6df061e0e621b63053c029719fd;
mem[737] = 144'h0b5ef3fbf2ff0302e9c6e736f5bc075c0053;
mem[738] = 144'hefa2e4e50243fb6f174617a9e3dffacf1902;
mem[739] = 144'h159f1f021abaf92f18eafd19edd7e5070753;
mem[740] = 144'heafee4dd0830f28f03da1619007106bb020c;
mem[741] = 144'hfb111073085d1348f2a8ea981e1bff00fc8c;
mem[742] = 144'hf22df8031adbf15307a8f26c1057ed170797;
mem[743] = 144'hf7c81df5e8a412dbe5b41ae5e8e0f2131973;
mem[744] = 144'h198ee05df625ffe0eff1126d07cbee16e15a;
mem[745] = 144'he75cfc70eee60c5404d803ec07010548f245;
mem[746] = 144'hf123ea53eb381a01eac30fae0164f99302b2;
mem[747] = 144'hee0a1fdb042d0d86ee17f31d1b75f21ef622;
mem[748] = 144'h171fe916e8f10a990f77e4a0f7980400f627;
mem[749] = 144'h1b5f195f002016d5e710fe3af233f6dcf09a;
mem[750] = 144'h1372e0e207ae0b69f93205821236f23d1f85;
mem[751] = 144'h1362e54d1839ebdcfe8b1af91fb318bc121a;
mem[752] = 144'h1670117bf4c0f6bfe85ef82e1f95f2be1a69;
mem[753] = 144'h0cf1135312c704d9149a04a41995e8dee15d;
mem[754] = 144'h108211faf3f1f11c1b440f4907cd0601ee5a;
mem[755] = 144'hef8d163507961fb1f64111470393f93505b0;
mem[756] = 144'h0159e7e111b1033befb6e6971ae0f421eae7;
mem[757] = 144'he0601dc3f9291c14f88d04e5e7921b0ae914;
mem[758] = 144'h1f080232e53ae83b0c03e87df05c1110e248;
mem[759] = 144'h1c99e50b168805820af0134ffa33feb9f440;
mem[760] = 144'hff4dff2cefc01c0d09ec0a68f9d9e1bd1e3c;
mem[761] = 144'h08f70e410bafe211e0c9e08ceb5cf5db14c1;
mem[762] = 144'he368e231f9b4f82efbededbe11ec16f51a3d;
mem[763] = 144'he7bc17b0f3a712ae0d1d03bb0286e2b2f079;
mem[764] = 144'hffa5e92ce72615bdebb6e26918401dceefaa;
mem[765] = 144'he6441585f921ea4af03aea3f02bbe1a5f7f4;
mem[766] = 144'h0deb03b3e7f2e7ea0cd306211622fbe61a3f;
mem[767] = 144'heacd0e48fd74fc5c1a000ec6e7a212f6e874;
mem[768] = 144'hf1b2e66b1ccae754fe4a1709e158febe1b86;
mem[769] = 144'h006df0f9e4a10086fe5f13ff1232fd331de4;
mem[770] = 144'hf323e85e0d5afe45ec3be69b0cbef1ba1301;
mem[771] = 144'he13f1e821a45fc220aac105de34714370777;
mem[772] = 144'h0b3817bf178d04c7e8361061edcae8a21dcc;
mem[773] = 144'h1e16e6130452e4fff3a70c3e089de8a1180a;
mem[774] = 144'h051610c40c8a1cbf10a8e2a00b9f1f9d165d;
mem[775] = 144'h0f91ec7f12751a78e1f8f834eb370bc90d6d;
mem[776] = 144'hf6fd13381ce1e057002ae59009820214e428;
mem[777] = 144'hfe2ef8d60e96f4af13530125e463153c1711;
mem[778] = 144'h12b8f0521beb1039ed280733e1d1e698e4bc;
mem[779] = 144'hea36e852e70efa9cf141e5cae7df1745fed6;
mem[780] = 144'h160212ba183f0d8af07c12f71685eee4e544;
mem[781] = 144'h1b73fd5304b70183f0e60eee12f21a0f15af;
mem[782] = 144'hfac915aaf090ec34f6da0b09f1d31078e265;
mem[783] = 144'hed7a06f3f9bc007af4240042e6d9f1410056;
mem[784] = 144'h083f0c0fe3b91d3d0554e211e12dfd81f297;
mem[785] = 144'h1568e167e907f2a2e36306b0ed4b13aafb79;
mem[786] = 144'hfacefd890593ea4be3391e2cf19905f116ee;
mem[787] = 144'h06e1f6121935e9b1fd161f83fab601ebef59;
mem[788] = 144'h179c0bdee1b1ed0d0712f48ee8b21b661c7d;
mem[789] = 144'h01f711ece5541cd1fa6506e3e970e93e0335;
mem[790] = 144'h1bfe0488ec131465ee8919bde29af4c7e8f4;
mem[791] = 144'he755102b0ba5102103b413c50111ecad1318;
mem[792] = 144'hee2b0d35ea961da3fa79147503e70dda0bdd;
mem[793] = 144'h200012a1e5de06231d50f0fc1ccd17220225;
mem[794] = 144'hec3f1091f2a6fc810cd9f545ef86faa8eb70;
mem[795] = 144'hf7a4ee7ee070e0421d54fe8002ab1c5b0932;
mem[796] = 144'hecb8145c1091067ae7e2e06be621f48510ec;
mem[797] = 144'hfe381be7e7aa0f1f0298e314ff4fe704e0a1;
mem[798] = 144'h0bfae6200500fa8e1fbc181f0045e759eb20;
mem[799] = 144'h099f04bdff4eef5e117ee8fe11c31ca6f708;
mem[800] = 144'h0139117efc17e06f02c9f1e1e998f3fdff84;
mem[801] = 144'heb60eb1f07fcf056e5f016c9e4f2fc7fe8d1;
mem[802] = 144'he392fc2cef4fea2b031a0f47fb010573fb56;
mem[803] = 144'h027bf1c0f61911ccfc9aecff0d8a1ca112a1;
mem[804] = 144'h107200c3076503890745ef3ffc481d4eff77;
mem[805] = 144'hf5afec0d000fef7ffcd41c54ed6df51b0563;
mem[806] = 144'hef46ea5e144be819ee581dbffd100f66eec4;
mem[807] = 144'hf4bc01f5f8df13cc1f58e253e196ea321e16;
mem[808] = 144'hee82eefa01c214ff10ec1f97ec76e0331a93;
mem[809] = 144'hf601090b04c7039e11b6fdec0b7ef0b709c6;
mem[810] = 144'hf9dc1aa2e9360c72f02ae6f20daf128c11b3;
mem[811] = 144'h0ccdfe3fe58c171a0d83e581190fe4c601cc;
mem[812] = 144'hfa3a16faf0c01cb5f9c3e31cee28e284f6b1;
mem[813] = 144'hee51e119e3161676f82c1d7ef479ed6500c3;
mem[814] = 144'hfd59e57f1f3812ceef03e42ee4f2034009c9;
mem[815] = 144'hebe7118ae18010e116060fddf3ff0ae51271;
mem[816] = 144'h1a0805bce664097fe4b6f813fa1e0dd5ff6e;
mem[817] = 144'hf195e4440179fcb1f02fea3cfb90f66de59c;
mem[818] = 144'he1fa06b8e41af12de09ce0e3f76ae7c805b0;
mem[819] = 144'hee7df4401fc50f6fe117f8071846f4440d29;
mem[820] = 144'h1efe0775ecb1edb4ef0915bcee371f50eab4;
mem[821] = 144'h05e1e09be582ede7eecd1079e235fd1f01f9;
mem[822] = 144'h1613ec94f4c30ecbe0f6fb2813021015f80a;
mem[823] = 144'h073319be17800e87f0fced1c12161801020a;
mem[824] = 144'hf007f9ee1fce1051f012ea6de548f8160ee7;
mem[825] = 144'heeb8e1b8ee36f09df573ee090eb8e24f1d91;
mem[826] = 144'he645f32e1a740fc6e565144cfbe8015608b0;
mem[827] = 144'h1904e7d60fd01ee0e036fda4fa3df2211b9a;
mem[828] = 144'h03080ab0efff101e06690d430fabe4b8f01a;
mem[829] = 144'h1f34e3d8ff12f44de5b105fdf779f7c810a0;
mem[830] = 144'h05fd10d818e11a25e609ed59034e1c2ee38f;
mem[831] = 144'h133ef5abe0201c5b1966e5881d5e13980b35;
mem[832] = 144'he2d4faf80815ec3d05f7f68de0d908e2f47a;
mem[833] = 144'h08641150f4391837ea770f320f9d14ae0b5e;
mem[834] = 144'hebf1e821e037107515040b77e542e508e5de;
mem[835] = 144'h1ae0f58918fae59c17210d5b067f05010f39;
mem[836] = 144'hee1215481758032516e3faf9ef1cee400d7f;
mem[837] = 144'h1918fa5cf021e7021ac5ed54119ce08d1704;
mem[838] = 144'hfcebe1f0133aef4e0576e9e104360f0eed00;
mem[839] = 144'hfec6ff03eb9b161bf5090b9d08d60971f9ab;
mem[840] = 144'h011a0d111a32101df0121a740e93ee5315b7;
mem[841] = 144'he48ee565e5abefa00f48196b0467f790f6f0;
mem[842] = 144'h1313e1521b2be9ace5f3e492ff6fe9c2e918;
mem[843] = 144'h16f1ed04e32efcf5f71e0439f73de3a0f0ea;
mem[844] = 144'hff101485171cf2711716fd7bfc39e9ce14eb;
mem[845] = 144'heca8000f079b032f0cec061c02330c5cf888;
mem[846] = 144'hf1ce06ed1081f8f810e9fd54172c048e0933;
mem[847] = 144'hfffbe048fb5ef96becf2e0ceef5817b80f71;
mem[848] = 144'h1be41ed8e9350ebb04a8e78ce01a10ae0d4c;
mem[849] = 144'hf9bd1ded10331e10fbc10de9eae913610b05;
mem[850] = 144'hf1560657ec1a06fd1a26ff12e477e20df009;
mem[851] = 144'h1be70314f749fe1b1c05ea77fdc2ec2de8dc;
mem[852] = 144'heb12e0ad1b68e477e7610a3df1a0f78d106f;
mem[853] = 144'hfd05e902eb1002801483072cf06efa100076;
mem[854] = 144'he3ffff701438e7250ee61f5306e00b2b0ab6;
mem[855] = 144'heb981e81ed9a076b1fe407b501f404f215cd;
mem[856] = 144'heb6df2e209b7eb84ffa706de015f1b5c1342;
mem[857] = 144'he1eb0472ec3ef5321f7fecc0ffadfe26142d;
mem[858] = 144'hf66b0be2eb4f0aae1f380805ebe9ea5e0811;
mem[859] = 144'hf3d0fe3eebe614d9e512f6f5e888ed4b0744;
mem[860] = 144'h16b71198e08aff92e4220ccc1757099af392;
mem[861] = 144'heec519581717ea46f7e7e437faeffdbcf133;
mem[862] = 144'h17fbe165e507e23216c3ecace4ddfe3ef71f;
mem[863] = 144'h1afd194809b20a0c073be93d0466e73413b4;
mem[864] = 144'hf3460f38edfafa7d10310a2ff427188de4ab;
mem[865] = 144'h0b6ef8e0074ae33ae08c02241044ebe9ec73;
mem[866] = 144'he446e881ff701de20d26e239e7cdeac30600;
mem[867] = 144'hff46f241121bf2befea4f4bc1430f91be05a;
mem[868] = 144'h1b0e016916391712187be24ae8d70da5feb6;
mem[869] = 144'h0d370281e268f0391d480de81272ebcb0f90;
mem[870] = 144'he4d9e77ef44aeed817c10cb6101e1f9fe804;
mem[871] = 144'hedcaeec01d9807440a9f1792e9070523eaa4;
mem[872] = 144'h09fc18d5e86af3b81ef2ee60014af7bbe6ca;
mem[873] = 144'heaff1bb01fb4188bec7c0aadf91bf5600b6e;
mem[874] = 144'h1a931eabe270e91c1f2d1214ef8cf47ce5fe;
mem[875] = 144'h0cf8105df585fb0df138089c19a2fe8b0e7c;
mem[876] = 144'h04fff06ef30df414104ce766e64af5aff1e3;
mem[877] = 144'h0da4ea4f064ef4f10752fa3ee666ef621a27;
mem[878] = 144'h16ddf7b8ee1e18e3f92f0a460f88f6ecf9b6;
mem[879] = 144'he9031a61e7d4f43c0fa8f6cbe0031890196d;
mem[880] = 144'hfe45e17119c1f1d3e5760867ef4719c7e1ea;
mem[881] = 144'h1ac01522090e0494e673f429f8effd5e0b6d;
mem[882] = 144'hf556e7620774117eef93e7530b62018b0151;
mem[883] = 144'h0ca61a9df503fa0a047813c7f49e1fec0f44;
mem[884] = 144'h1988f891e27ced56f8e40f69eb4ae1df1589;
mem[885] = 144'h1a5d035317f81578150f166d06c1178c16be;
mem[886] = 144'h1265036fed031451e4f70bc20b1dfc271597;
mem[887] = 144'heb3f0dcdfbc3e09eedecfd16f145f803fe5a;
mem[888] = 144'he987e4030e5c1bf10e940c34e18318630dc2;
mem[889] = 144'hee14e943e037fd7eebeaedebe4af0ca4ef79;
mem[890] = 144'hec6bf022f8970b141892e0d2e460f5e6119d;
mem[891] = 144'h14730c65e9a2fe35f2f5fa27e53f0199ed42;
mem[892] = 144'h1604fe8b04b8e89e031c17711233e41c1081;
mem[893] = 144'h0307ee8401be074ef4c8120cf5c6eb111d33;
mem[894] = 144'h066be2a3f2f61456ecdaf8f6193bfd1ffe5a;
mem[895] = 144'heb80faa81932e4591032f383153511e1f7fa;
mem[896] = 144'he72bf03916c4ea37f68c03e3f6f6f850f8d2;
mem[897] = 144'hfc9909940d49ee6c146312f0e33b10b6facf;
mem[898] = 144'he331fc38e7d904aa05b6e4e7ee0315d71a7d;
mem[899] = 144'h010f0aecea07fb891f8aee03f816f5ff13e4;
mem[900] = 144'hf824e3c301beef46f3301fd8f7d4062b1593;
mem[901] = 144'he71b0c3de3ace64eef16ff72e1d10308e74e;
mem[902] = 144'he6dcf79eea56ec9bfbaef95b0ed10d0e0cfb;
mem[903] = 144'h1f2d0739061d040a045f19b51dcb10d5eabf;
mem[904] = 144'hfaac07e00888f1a3e8d20cf7fdace6981e84;
mem[905] = 144'hf7dd0787f445e314fcd80a3df76cf32ee0a5;
mem[906] = 144'h0363f7f610b20a8c10b0f00a1ae3fa2712a4;
mem[907] = 144'h0726e65ee274ec8ef39209771242ed90f96c;
mem[908] = 144'hfbd8027d1cc11d15fe23143c0bce1c001c08;
mem[909] = 144'h017d1d560ed01b5e02b216a7e5adf46e1429;
mem[910] = 144'hf48fec1c041b0d08ef300409180310e30125;
mem[911] = 144'h1bc013a70a35e0f5006e0b0cec2909db14a0;
mem[912] = 144'h00e5f85deae1f7b7e5010b3310471dfdf846;
mem[913] = 144'h0ee40ee816dded8bf91c04f7fc89f6771c44;
mem[914] = 144'he66df122e874fcce1c0d06d2ef01f38c0a5b;
mem[915] = 144'hf23c12430f5117c1f9d9f502e8cd1a240422;
mem[916] = 144'he8c80db7f749f85b1030f8961f27f6400480;
mem[917] = 144'hed691787fd6c12c2067116c9194b1722fb6a;
mem[918] = 144'h1f3bfa7b1a54183013561eecf7411782f2d2;
mem[919] = 144'h00260066104316a1f64be7e900a9e317ed95;
mem[920] = 144'h109405be130116d607781c4bffaee131e5cd;
mem[921] = 144'h1872f6df0cb30818e1daf1751087efb4e75a;
mem[922] = 144'he9af10240068e165e77b1e28f191f87df1b3;
mem[923] = 144'hf2daf80ff328f1e6e73b076616bfeb601485;
mem[924] = 144'hf504f40e042c10a2fe70099a0afbf3410d97;
mem[925] = 144'h09aff0d1e42f081d1118f5aa14b3f09bfaa2;
mem[926] = 144'heac3e06518831f1be01b0274032819f71dbe;
mem[927] = 144'hfc7dfec1fc3f13c013b01844ec5aea2b1171;
mem[928] = 144'h1e6104b10eb2e51b184df23419fef370e7da;
mem[929] = 144'hf261faebf5c305cde6e9ffe9e085e579136e;
mem[930] = 144'he4911c6af41bf25f194feef5e09aec35fff6;
mem[931] = 144'he09aebb6086e0d43ee11fd9109d40ca6e390;
mem[932] = 144'he91b11cde47df264f0f901df16f7fc7b121e;
mem[933] = 144'hfed6e0f906d703ec02b00c31f763e386f28d;
mem[934] = 144'hfff8f38b0d4410ab00e919dd194be41b1031;
mem[935] = 144'h1fbf0ae60c4efcefe2e8ecd9ff73f87afc7e;
mem[936] = 144'hf07c12890fe2ff630f8ee27eef97e1cc1519;
mem[937] = 144'he9df1452f0571be3f4c8fbbbeba00ffd01d2;
mem[938] = 144'hed65f8a5ffe7f3781a510b1b1f4e011f04ca;
mem[939] = 144'h0c6ffbdce704eef41ccd19d6027a0f2f0737;
mem[940] = 144'hf8eaf63b0299e41dee08070ff4901853ea6d;
mem[941] = 144'hf0c608aee16b1fecfaa612ae088b06670140;
mem[942] = 144'h114e15eaf1cd11e3fcab07870fe501c3e893;
mem[943] = 144'hf57de3d70405eeda1a87fea4e9821bd90537;
mem[944] = 144'h0e1eefa21b6ee962e983e8c5f00f12fc03b7;
mem[945] = 144'h100a093b1a52022f1d1b00fbee97f9f7137a;
mem[946] = 144'h19d90110e59f101e06c9e90f0e7ce41e0893;
mem[947] = 144'hf2bfe9040664e0ea1774f68be1a0e1e7f4ad;
mem[948] = 144'he06f0ddeefe3100901a312300efae95afe73;
mem[949] = 144'h12800b41f675e0011164e728fa8000681745;
mem[950] = 144'h0f68f7a9e7b917def9a9e9601e21ebd8157b;
mem[951] = 144'hee831abbfc69f58a19761867f1e20483ff4a;
mem[952] = 144'hefb20628e230e869f5d2e738156ee9f2f1e2;
mem[953] = 144'h04a10461f410087bf4d51eae00ecfae4fc7a;
mem[954] = 144'h09e1f6d30a22e7eafbc2f32919d41b8a1b37;
mem[955] = 144'h0b1befa31b2df98611a31dcaf9b002a70036;
mem[956] = 144'hf42d0662fd89fc4d09e51f96fa89f3c1097f;
mem[957] = 144'hfee608aeeb69e606f10818c4ff5b18071878;
mem[958] = 144'he1be1e45e6751cbfe55feb61e52bf383127c;
mem[959] = 144'hed96f6b8006b0c18ed10e7f8e35fefbbfe91;
mem[960] = 144'he3431869f21814971548f3ea015dffe30de2;
mem[961] = 144'hfa5df4fe08370ba9e0b1fff9fbfc01dd08d8;
mem[962] = 144'hf3f4fc7ffa2ae60a12b601ee03e81c8be587;
mem[963] = 144'h0aa7e391ef65e1930c19e4b5eef4fecd1bc0;
mem[964] = 144'h13b5e7ace3c8f469eeacea6105bfeb4f11c5;
mem[965] = 144'hfc351f1cfc8f021f181e1c061b23e94fe445;
mem[966] = 144'hf693f2ab08fce1b9fdcdfbc9e0b9e05bf163;
mem[967] = 144'h1faaea980768e572efe5f4ebf4830c521e42;
mem[968] = 144'h11471639002e06f6f3c409011ba30931e324;
mem[969] = 144'h07671f20f2d10daf0494e649142d0ef0ef1c;
mem[970] = 144'h1d8e1294ea0505a214e7049b0a89e201f5d5;
mem[971] = 144'hefed069f1273e29e0b94fb8affe6e27502cb;
mem[972] = 144'hecbb1a69f2b212cc071ae1b0e081124ef5ed;
mem[973] = 144'hfd86fef3fee1e273eda317711fb5e8fdeb2d;
mem[974] = 144'hed0cf96bf10ae0c01ab1f4fcf18600c4f59d;
mem[975] = 144'hfb34eebfe2e0e92518de01cbf19708910c03;
mem[976] = 144'h105709de10ddfddbf415e671f7b80119f9a1;
mem[977] = 144'he182e1170a2511b4ff53ee3c133a11390473;
mem[978] = 144'h05e0f3c0f212e6d615841b8a0354efaae29d;
mem[979] = 144'he9ed0793f212ef2beaf900551ea40b521694;
mem[980] = 144'h14caf4b6eecee6dfe39c19b1ef49054e1958;
mem[981] = 144'heaec1f1a1303ed95f79fe074fd23fc0f0736;
mem[982] = 144'he4ad17e9e988ef31f797fa1302e7175e0196;
mem[983] = 144'h1434eeeceab31946e236ecb81b57046b095e;
mem[984] = 144'h0101ea28f80e0e51ee6811c31f26125f02d5;
mem[985] = 144'hf99109cc04f7e246fa181151fea1fdc3126b;
mem[986] = 144'h0ff110970d4b0744e5c6f03e06f302ae0468;
mem[987] = 144'hf20a19cde5caebdc01be1e64f83fe885ff85;
mem[988] = 144'hfb90e95902cf1a5d1edf1215e07de459f2c1;
mem[989] = 144'heebc0710e704e17bfdde0c3b18ab02480dda;
mem[990] = 144'hef5e0b16f862e691fc1ce18b0eeb1aa9fe06;
mem[991] = 144'he4aae3ad1e4913ca1e2dea7e1fa7f0cf1ceb;
mem[992] = 144'h064113b0092f1a8bfca3f6621946ebe21f9c;
mem[993] = 144'hef07e68f17c40e42eb24f97c0fcb026dfea8;
mem[994] = 144'hf824fe0708590f0803d907710f7b07ee100d;
mem[995] = 144'hee6f05c1131d064ae091f1831c5af9c10bf4;
mem[996] = 144'h1a8f17701bde139814faf3dcef84fad31d36;
mem[997] = 144'h17e0fcc41407058a1467ea6a1d0ffca2f629;
mem[998] = 144'h149f0927e537fa4103f51ba30d3f03e4e0a4;
mem[999] = 144'hea8e12220985fc76e8c7f0d313cffa411d95;
mem[1000] = 144'h1c471ce7192a0528eb49e2bd09b5f6ee12df;
mem[1001] = 144'he913ecb5fb45fd510aa11dfef642e655038d;
mem[1002] = 144'h1eade45d0437129cf2f9e391044d003b0fa7;
mem[1003] = 144'h13ed015f17b3ea0e123b013a1dabe4dd15cc;
mem[1004] = 144'h1809088fe8581688e5390a3c0528f91e0b63;
mem[1005] = 144'h092c1c290a00eed0078bf8adea2c1dbcf76e;
mem[1006] = 144'hfbf80de6ea2dee30f82c1c6e06cd11a201c8;
mem[1007] = 144'h11e60b760d6ef25f00a90e6af3bafffe1a63;
mem[1008] = 144'h0f5ff6c11932eb370bc5ff9e17711552172d;
mem[1009] = 144'he3c8108a18aa03e31af0f1f1ea991beb1bde;
mem[1010] = 144'h1ce611e2ee10f6b2e00b0c2714c7ed3af4b8;
mem[1011] = 144'h182bf80105901b47ead204541ecae9ddeab4;
mem[1012] = 144'hf6550b3613a1f022e7690b7ae136f35ee867;
mem[1013] = 144'he1b9f634f34dfd930d63085aeca4f45cf12f;
mem[1014] = 144'hef7c10150fabfa57035af9331b74e5b80f81;
mem[1015] = 144'h12caf14befdd1930f002029d1531f261116b;
mem[1016] = 144'hfeb70a75ebb40a91e2130bc8efadfce9029f;
mem[1017] = 144'h174de57201d7f282fb72e77412a204e51f72;
mem[1018] = 144'h0715f2ab15670d8cf5d0ec25ef46f924141d;
mem[1019] = 144'hf8661a2a01abe51b00e304b8f0d41801fb5d;
mem[1020] = 144'h062d17eb1e35e981071219bde2bd1078fb31;
mem[1021] = 144'hf4ba0a0218ddedb600a4eed7e4fae146112b;
mem[1022] = 144'he8f019a2ed22ed050bfb0b53ee3910991774;
mem[1023] = 144'h08890aaef7b8e368102f1630ff4d143013ad;
mem[1024] = 144'heb2eecb715cf120f17a8f50cfa88e09b0f58;
mem[1025] = 144'hf8e30151f7240b0fe2a412fa0bb91ae31189;
mem[1026] = 144'h0f88ead809e1052bf019ef07f937ef81e447;
mem[1027] = 144'h06c6e173f352f567ed37e1c5e44b03eb0b81;
mem[1028] = 144'hfd3aef51e270004002affd63143efd1e0817;
mem[1029] = 144'hf7211ebfefb20c140c9ced1212bc1b5a0487;
mem[1030] = 144'he3a41466ec59ef36ebb5138ce233fb251deb;
mem[1031] = 144'hf83a0e1f010201c1f841e4bc1b8a0e0619ec;
mem[1032] = 144'hf589182ae76a1769e836fb4aff81f8b1ed6c;
mem[1033] = 144'h0ee2e8221ada1dc71c5c0c38e691fcc4ff32;
mem[1034] = 144'h0586162b12d21c42f082f90cf3f3e0a519f5;
mem[1035] = 144'hf75e15f9f8a9f1a5ed1911320133163405de;
mem[1036] = 144'h12e00269e4ec0e7011300e45e650f7f51863;
mem[1037] = 144'h0d88e563ec15f69bf1bb10d008d50c5a0892;
mem[1038] = 144'hfac8f426e7a20d8909d5f38c1ffc1396109b;
mem[1039] = 144'hfdf2e09cff5d112406a90298ed061aca0da2;
mem[1040] = 144'h1d18fac21443e32bf2371cf40b680a69efbe;
mem[1041] = 144'hfd3815431efaf58914e7f678ec7008730f76;
mem[1042] = 144'h18c3e168ec5ef320fba3ed3ae8b10f8c1b12;
mem[1043] = 144'h0963ea30f2f1fc5a19b30746ec7d1cc1e516;
mem[1044] = 144'h0952e1d31df6e28d07fb0a820da1f9d90ff9;
mem[1045] = 144'h178dff4bf911efb3ef470c1115560e46e885;
mem[1046] = 144'he39e13d7e00c180e0b2fdfc21a86e3421e78;
mem[1047] = 144'h00140529043dfd001c420ce910bf129be194;
mem[1048] = 144'h0f7be779f9c0ffd813b31149089d1969f331;
mem[1049] = 144'h0d771f0de26dfac5ff5508a615d40b4df931;
mem[1050] = 144'h128de18ae19efed911391b24fc031eba1892;
mem[1051] = 144'hedb3f0abffa9e50efef4e2c6fccdfffa1c97;
mem[1052] = 144'he28f10711afced52f2a3e4f2e874fbc3fcd0;
mem[1053] = 144'hfaa1fdd4e5e70102f7c9f0caee4004de152a;
mem[1054] = 144'hecd40f05e0601154f0f2f30c1e3a13361083;
mem[1055] = 144'heceff5e91acc0c070f8efcec04eeea66f2d5;
mem[1056] = 144'he6e50b5dfb34f085eed5e1e30a4f0a2f019d;
mem[1057] = 144'hed40040de4951e6c10f6ea121720f701efe7;
mem[1058] = 144'h06550d5de60f0dadfb90e265ec8ae9fee37c;
mem[1059] = 144'he46e006fee6ae6580d63fb1dfb1a1d6503e8;
mem[1060] = 144'h0b1bf0e31b8607f3e0060bb51197191bec37;
mem[1061] = 144'h0f31f43fea921bffe8c0034d1163087ee8ae;
mem[1062] = 144'h0d70f8f2e162e5b40926017604fbece50a77;
mem[1063] = 144'hec06193e0e30e0e8e23e08e40d8418481ba1;
mem[1064] = 144'h073c10820b9af293e977f71de3961c54061b;
mem[1065] = 144'hf0081da2fb72e2f60f98f53607fff25212dd;
mem[1066] = 144'hf836101efca402d90107ed3dfe0b197812d3;
mem[1067] = 144'hf35d1c07ef770de0e607e387ea62174df4a6;
mem[1068] = 144'h1822fee00b3d1e72e0e3faf0092cea6c0f8a;
mem[1069] = 144'h1d14f199fba71b5814a1e01e1b14e86012fc;
mem[1070] = 144'h124fee19e3f7e7cd0457e49610c10293171f;
mem[1071] = 144'he2f51c810143ff23e3c3013b1211ff8112a7;
mem[1072] = 144'hebeae9c5fbf20e3402920ff90f10135b0de4;
mem[1073] = 144'h028e078df3f817b1f1b1f167e463fc22f41b;
mem[1074] = 144'h0c2306bb1ac6f71218040a750e1914afe459;
mem[1075] = 144'hedfd126100590dc5e872094d025f1f5bfd61;
mem[1076] = 144'h1e750fe8e2f0f8ccea79ef82f2eefaebfc67;
mem[1077] = 144'h09fcf86910140bfaf2e4121bf8bc1c881bd8;
mem[1078] = 144'hfb5ae2d5f9be0a9d143e0d87e8fde93dfadd;
mem[1079] = 144'h0af3073cf533f124f8340aaae0c00acbef63;
mem[1080] = 144'h07b0ff9510061fe11e5becb6e586ee260b59;
mem[1081] = 144'h1cc717e4e71407a7ea4e08c6f69a0e941eca;
mem[1082] = 144'h1251096bf2f7fe0df1fde3c1026d0eaf1dbc;
mem[1083] = 144'h0c98efc704faeaade8edfae901a40029e80c;
mem[1084] = 144'hed0a033af81e194ce7961a2b10ce1e44e0a3;
mem[1085] = 144'hfa9704b4ee06eb751d25f46d03ac1bf9fcad;
mem[1086] = 144'hfc78f8fef06b02480a96102deffcf56c146a;
mem[1087] = 144'hfbadef56086619750c6ceb3b07c21fd4eebe;
mem[1088] = 144'h16fd094e1680f2c6f8501f6af9ecfd87144a;
mem[1089] = 144'hf74906aa0330150b161ae79b1e23fe92f655;
mem[1090] = 144'h02b701eef95fe8341a061e850d8f0645e4b7;
mem[1091] = 144'hfbd6f34eec2e0839008b0e0d1d44edbce2db;
mem[1092] = 144'hff5effb9048bf24ae264ece5f89ae97a1e98;
mem[1093] = 144'h080505b41df30b2cf5ea04d808d408ea0e91;
mem[1094] = 144'h0001094cee150330f1ea0107e51e0adf0c56;
mem[1095] = 144'hf5e6fcd2f345f7fdf59411071da01d20128f;
mem[1096] = 144'h02e2e6dae05607cde253fc821eafe289ed40;
mem[1097] = 144'he3fcf9fe1dbb1326fa6ef25611c5eb840c52;
mem[1098] = 144'h0221e66feb5001b41165e30406901e0ee1d3;
mem[1099] = 144'h096b12190581033c013008a50fd014e61d29;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule