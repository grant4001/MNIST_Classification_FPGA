`timescale 1ns/1ns

module wt_fc1_mem0 #(parameter ADDR_WIDTH = 10, DATA_WIDTH = 144, DEPTH = 1024) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'hf4c6f700f1a2fb76fa14051a0c18fde80d31;
mem[1] = 144'h0be00176fbe8fe92fff2f2820230f823fd97;
mem[2] = 144'h0663072af5fdf921f5930daaf9adfeeb050e;
mem[3] = 144'h01b40e610ed2ff8e04440956f0ac091c091a;
mem[4] = 144'h008204d2fbd4f3a3f159f2e1f72d0889fed2;
mem[5] = 144'hf202f01f0c2f03daf6cb0f9f0722f70df86e;
mem[6] = 144'h01060ec0fd53fe000f21fb52fba703650b3a;
mem[7] = 144'h0f290243f320f744f73a0c9cf90bfbcd02bf;
mem[8] = 144'h08acf69f067afde10acef002f438f1fa0c83;
mem[9] = 144'hf1500dfb06080eaafbda0ebf0aa508d5f701;
mem[10] = 144'hfc1df8040afbf515fe38099c017afb250526;
mem[11] = 144'hf69df09dfae0f7610dacffb3fe1eefc00d3a;
mem[12] = 144'hf506f51602c3fd010b92f695f7460f6eff1e;
mem[13] = 144'h00c30794f4c707a40595f50b0e1c0423f482;
mem[14] = 144'h0d5efd2a07b3fdb80fae0943f8d00dea05e4;
mem[15] = 144'hf90103640c59f00ef487fcf9fc3bfa1bf5c9;
mem[16] = 144'h064af2aaf850f3fe0fce032e01d9fa4303a7;
mem[17] = 144'hf4910c19008b08d8078e0787f631f1bb04f4;
mem[18] = 144'hfb41fd03f57a03ed0e6bf30808a50a9cf5aa;
mem[19] = 144'h0f760eb3f8fffac70cea0f1005800e61f0bf;
mem[20] = 144'h08b200a2f2130576f8fcf67206a5fb2306ab;
mem[21] = 144'hf079f9f40d52015f0d61037bf0e8f4740d2c;
mem[22] = 144'hfcb6fd26f3c0fac2f0eaf3def09b01680b0b;
mem[23] = 144'h00f4fb0bf7d7f6510358f52f0b80f693fff9;
mem[24] = 144'h045cffbb07490025fe980007027cfc39f2f4;
mem[25] = 144'hfc69fa7306c305c00b0509f8f045fe7c0eef;
mem[26] = 144'hf80ef144f6a0f623f8800c0f068d002df318;
mem[27] = 144'h0fa5f66704a3087600a1fcedff41f9990524;
mem[28] = 144'hf6ad0bc70e31091cf230f37e0b1b0d7e0ecc;
mem[29] = 144'h0fd1f8c8fd8ff090f870f6baf15c0c7c0afb;
mem[30] = 144'hf618f3d0f7e7f8befcda0747fa160510fe81;
mem[31] = 144'h02ce0f600f3b078bf038f65907aaf8a4fd5c;
mem[32] = 144'hf41af1c201bd02280de2f73e07f3f220f009;
mem[33] = 144'hf66a0f7df2b509c1f3670a47067d049f01d0;
mem[34] = 144'hff95f574051ef4f50ebdfd48ff6d0a520122;
mem[35] = 144'h0117f72df24307a5092f0779051b073a0e76;
mem[36] = 144'hfbf7f22f05b006edea39e252f84dfe58fcaf;
mem[37] = 144'hfe9a08f20229ff710764ecb1f1280285f9b0;
mem[38] = 144'h02fc0b6cf86afa2ef3f6f8200d500cfb0907;
mem[39] = 144'hfdbffd3a02bcf53b01b8f6de05d7edf4f2ff;
mem[40] = 144'hec87fb9feb2eec72f503fd5efb2beef5dedb;
mem[41] = 144'hfff10b1eff4af6d2027800f808d803afee22;
mem[42] = 144'hfe8e09d001cafa30f6b4f9c90c9cee45ef08;
mem[43] = 144'hfe0af901029cff5204880d940a12f11b021b;
mem[44] = 144'hfb8f00acfbd3fdac070401dbf7e6fb0505d9;
mem[45] = 144'h07950d13ff9d047400adfff907c8f7c60c2a;
mem[46] = 144'h094504fa0ae9f6c50fd804ea0cea00360ac3;
mem[47] = 144'hff510d8c095a0b3ef35cf7400b32f028faf0;
mem[48] = 144'h0e410763fbf0f9880e8806cc0bd9f0dd01ba;
mem[49] = 144'h03d4f0300c8903d20c16fae804aef8410640;
mem[50] = 144'hf8c4efe4fbce0d75f7f6fa5002e0ff900bb0;
mem[51] = 144'h0476f7a6f364057d0295f89efb42f03af6a9;
mem[52] = 144'hf0b1fec104b4f1e3f7ee020500d1ef33feac;
mem[53] = 144'hf5c4f1faf91207bf0a8d0bbb08e0f5850da0;
mem[54] = 144'hfacc0cf3f13df30ef0f0fc7cf65cf59100f3;
mem[55] = 144'hf76405660277002dff75fa51eeae0342f908;
mem[56] = 144'hf601f352f9ad0620f4e0f601fd3eeda6f3a0;
mem[57] = 144'h09700d3a02f0f169fe32f05903830676f7f3;
mem[58] = 144'hf99ef6dd081cfb2af6280624f8e7fcaffb35;
mem[59] = 144'hf6a1f5f6fcb7f1b30e6508f6fe33fac10a1e;
mem[60] = 144'hef5df5c3f8f00a7cfdb8f517049cfc6ff6bf;
mem[61] = 144'h0b860793f005f69b027efe4b050aff430ab4;
mem[62] = 144'hf8c001a3ff2500600bf70f3c0a1b0d160201;
mem[63] = 144'hfb62f802fc5f04c5f17208fdf98800b80cc0;
mem[64] = 144'h0c4b08f8f4d7fa1e048d07190a520707f30e;
mem[65] = 144'h08bffac6f60dfb290098f428fa7505e50378;
mem[66] = 144'hf7d90be50bd405a8f8f50b120494087cf2d5;
mem[67] = 144'hfa86fb21f430fcfb0a690694fc7cf40d06cb;
mem[68] = 144'h0e2b022cfd9deec2f096ff8bfdc8f7d5ee57;
mem[69] = 144'h083207b10ad0fcdcf6470693f734fe33ecae;
mem[70] = 144'hf5f508c9f0450020f6d50f1ef18e08d90ee0;
mem[71] = 144'h09e5f1f4f1a9eb8ee93ff574059c030509eb;
mem[72] = 144'hfb31fccdf94ff6a2f4aaeeac0230e73def5f;
mem[73] = 144'hfeb3055c0849f937f33505e4098af70df4c8;
mem[74] = 144'hf802feeef911f73ef5f50d280902fd3cfb71;
mem[75] = 144'h0d4f012ff821f5240a3404f7f742f546f1f0;
mem[76] = 144'h01b2090605caf5de0d4d099309def26502e2;
mem[77] = 144'h090d0967f7b00cb90d0ff00b0b54f0bc00f7;
mem[78] = 144'h0bc8fd7b0eacfbea04a7f80b0acbfa89f790;
mem[79] = 144'h0e300d3c0771f2ac0795fc7bf5af08cd0a97;
mem[80] = 144'h00760740f6b5f1a80735fb03f41c004e07a5;
mem[81] = 144'hf7e40111fc230c40f022054e00aff41bffc8;
mem[82] = 144'h0863fd07fed10a900ad10e55f2a101a3047d;
mem[83] = 144'h0f650bc500c409a5f4a1f2e700cb0733f060;
mem[84] = 144'h0016fa0af1fdfbd4fc7bf300f1c0f85cf129;
mem[85] = 144'h012c03070141f11cf8e3ffc60e61f03200a9;
mem[86] = 144'hf023fad7034af15af453fa9c013efbe1f788;
mem[87] = 144'hef3b096204eaf097ff67fd65088309e0fa84;
mem[88] = 144'h08bcf812f344ee3bf70efdf3fd5601fe0309;
mem[89] = 144'hf5a6f229edcc0a28f15f0659ffca09090133;
mem[90] = 144'hf5030c40ed70f034fbf10c77f166fdd107e1;
mem[91] = 144'hf37bfef0f44b0fb9f8c60ca5ff1bf8baf548;
mem[92] = 144'hf4930cb100caf607fe32fd1d02190ccaf456;
mem[93] = 144'h0761fa6305760bc80b44044d07a70a9d0096;
mem[94] = 144'hf406fedbfc83f3150292fe98fdcf0288f238;
mem[95] = 144'hf417f75efc2c07ad051e0bcb0318f7ef08f2;
mem[96] = 144'h05b7080008850ba6fa99f107f5f10da10b83;
mem[97] = 144'hfbce07d404e9f7d5f5160a83f0b800ac0df8;
mem[98] = 144'h029202b8fcc9ffe0099d0755066708810c48;
mem[99] = 144'h0c460e73fe9c09a4f9df0ce0f0fbf2840aa5;
mem[100] = 144'h0ab50aea035d0041f0a6f8ba041af532ffc7;
mem[101] = 144'hf96bf1ed0a0304f9ff66073001db0d18f088;
mem[102] = 144'hf430f2100dd0005f083d01befd8a084d079e;
mem[103] = 144'hf553f32004ab03c50973fea9094703d0069c;
mem[104] = 144'h04a9fa5ff5def638056af1c501020c3f09cc;
mem[105] = 144'h021d08e0efb70acaf005fadc06a20fb3019b;
mem[106] = 144'hff13ef19fe18f71c0861032b08f7fc9ef81f;
mem[107] = 144'hffabfafd06ae092ff49604880b68f439f5f6;
mem[108] = 144'hff57f814f7c5ffcaf05e0646f11f02a8efc7;
mem[109] = 144'hf9dcf2200d390362fdbff460f74f07b5ff68;
mem[110] = 144'hf93e0b8cf6f5fe37f3f6f249f87cfb350cac;
mem[111] = 144'hff54fda608c60969f259f27e0b6a0e9504ab;
mem[112] = 144'h0f380dea023afd9000550ae8f4b20e26f778;
mem[113] = 144'hfade0ead07c2f19ef82b0576f099f0e602b3;
mem[114] = 144'h010cfe2bf4590e48fbbf05e2f912f6aff76d;
mem[115] = 144'hf35f032cf76b08f8ff9d0867f6610c8e0620;
mem[116] = 144'h0bcaee27ea2ff279eb4df7460682f798fa8c;
mem[117] = 144'hff750c73f1ab072a0ada027cf72bf70ef3ec;
mem[118] = 144'h00e607a00694f101f15f0878002bf565f935;
mem[119] = 144'h03bc02a70335fab9eecc0b1501af06d6f215;
mem[120] = 144'h0de3f97bec0be476028e0396f276006aea18;
mem[121] = 144'hfde70db7ee4bf493f798f307f44308eff7e2;
mem[122] = 144'hff08f9e303e8054eff84f39ef9c1fb51fdd9;
mem[123] = 144'hf1a0f636fe1bffa10a96fd0903fbf7a6ff2d;
mem[124] = 144'h001afea70069f07af202f4b6ff30f919093f;
mem[125] = 144'h04bff999fd03f1f907eaf1150b1a090ced41;
mem[126] = 144'h06b50e3504600d3d0d6f0d6b08810643f3b7;
mem[127] = 144'h048b0c660bb808c8fa34f28cfcdbf90c0c76;
mem[128] = 144'hf402fedcf494f279f8bd08a5f0e7fd16f451;
mem[129] = 144'hfe97062ff5760731f133f473098bf3380468;
mem[130] = 144'h0fb10ca9fac90afcfb9c0486f773f37102c2;
mem[131] = 144'h03d9f8e6058bfff8fc83f4d8fd9708a7f368;
mem[132] = 144'h05dfff830ee0f2a1fa4cf5f30b96045b0d1a;
mem[133] = 144'hfd27f67f0d30fc02010bfd6dfb2f0439ff6f;
mem[134] = 144'hf4f802faf177fc25f6ab01980c950c2df091;
mem[135] = 144'hfe960c0404eff515f300ff65fc0bf50ef31e;
mem[136] = 144'hfc8eff0cf7cc048604d30c3cf4a3ff3705cb;
mem[137] = 144'hf43dfcc4fd66f99ffc9cf7990e80f4aaf41a;
mem[138] = 144'hf95d0c630dbf071cf471f46b08c6f53ff741;
mem[139] = 144'hfb6afbfa0aff07a2023df8e80c9bfb8cf9a2;
mem[140] = 144'h0899fd9a0c28fd35f6bbf641004101abf50b;
mem[141] = 144'hf07af005081109150180f01cf52dff45f775;
mem[142] = 144'h085cf2a3fe60fb38f9f70fe3041b07000151;
mem[143] = 144'h0b3cfa99fa7808c3facdf82704210b1ef02f;
mem[144] = 144'h08120918065b0cb706cf0037f049fb9b084a;
mem[145] = 144'hf577f8b50070086605adfc02f371fee50650;
mem[146] = 144'h089af5b8fe08f39bf8adfa1afa110616ff91;
mem[147] = 144'h0bdef2bef389f48bf888fd25f4640f510afe;
mem[148] = 144'h00890cb20473fca9037105adf07a09ea032b;
mem[149] = 144'h00c200baf49cef880527f74cff0d0e52f500;
mem[150] = 144'hfd9c01cf0b4d027e0f05f918f212fdeff88d;
mem[151] = 144'h09bf0d95058bfa58fb83fddbf5bef198f7e1;
mem[152] = 144'h01b203dd06930e990f040d17fe9a0e5bf3bf;
mem[153] = 144'hf62cf31508e2f5b801b0fb40f02001a3053b;
mem[154] = 144'h09cd0b4ff65cf32d03f7fb1bf189fe840a66;
mem[155] = 144'hf739f1b1f0fdf476fd43f03c079e0046fbf5;
mem[156] = 144'hfbec0035fa0d096308acf741f424f6ba087d;
mem[157] = 144'hfb420c37020d0de6f692f0190a6e07b0f26e;
mem[158] = 144'h06ad00ddf59502620dbafc9ff6ba07c8f129;
mem[159] = 144'h0dd20013f00ff58dffbef101ffd8fa00f8e0;
mem[160] = 144'h0a77fd83fcd4f8fb08e5069f0315f739fa0b;
mem[161] = 144'h07dc0e6f0fd90cbff0e605b5060a06bd0b82;
mem[162] = 144'h02c1f2f9f4630df2f84d076df8ff07a00ad0;
mem[163] = 144'h02d7f675f80302ac0c6b0e8e0f9dfa130a1e;
mem[164] = 144'hfe24ff9ef34f03e1078501bbf4d50689ffc0;
mem[165] = 144'h0efcf08ff401f045f379f68df8cf00dd032d;
mem[166] = 144'h0d7d05e2f19c0df1f89aff72f2770c990fb2;
mem[167] = 144'h0e7efd3bef1ef2fc0bc800f9fae2fe3f0dcd;
mem[168] = 144'hf8f3fec108d804880e8b0e4806e1f51703d3;
mem[169] = 144'hf58401110e00fc3d0f27fa88f22cf8f6f76a;
mem[170] = 144'h073009dff794fcc20874f2550266fca80b65;
mem[171] = 144'h0919f008f999f1500be9f6c1fbf3fc5903cc;
mem[172] = 144'hf36d0f3ef8c50dadf760f04607d4f517f2aa;
mem[173] = 144'h0210fb81f3e6f25b0362f8a3f050f9aa09a2;
mem[174] = 144'h0632f264f510f403fe1df0c8fec20357028a;
mem[175] = 144'h0abe0388f4c8fe2ef297f254f8f70eccefe9;
mem[176] = 144'h09010e31febe039df2960950037cfe2df802;
mem[177] = 144'hf3220d0506900872ffed007c08cd0335fc1a;
mem[178] = 144'h094df1c70f4506040fd2f50bf801fca3f19d;
mem[179] = 144'h087f07ca02d20d03f9abf5fc0b1e075fefdc;
mem[180] = 144'hfc27ff5cf24af375fdd6014500bef58600d0;
mem[181] = 144'hf22a024cf865f7f10333fa23096ff0d6ffec;
mem[182] = 144'h0a73040009fbf083fc510541f640fb59fc02;
mem[183] = 144'h0b10044809e706490493057c01ccfad60e58;
mem[184] = 144'hf758ff8e081c00fafe000b46077002edf861;
mem[185] = 144'h012603b9fde90eb0f848f732014e0b82f116;
mem[186] = 144'hf571fe9cf8570f04fe71ffd101860fc7025e;
mem[187] = 144'hfc71f6a7f285f4c9f078fe95049dfd9af465;
mem[188] = 144'h06150c64f1dc0e260d2dfde70d50f1fff75b;
mem[189] = 144'h0627f4ab0809f39bf3ba06e2f0d9f859f70a;
mem[190] = 144'h0cca0a0a03c3f3f805d40bec07ddf49e04e6;
mem[191] = 144'h0062faba06dc09ee0141fae9018a0372f45d;
mem[192] = 144'hf619efd90677051ff706fa900cbaf6bbf58a;
mem[193] = 144'h0c7dfe87f2710e2fff470f3b0939f656068c;
mem[194] = 144'h0161f145fe03f9d0f17a0852f30ffabd079f;
mem[195] = 144'h07e405b3faddf9080a34f8930cea08c603a6;
mem[196] = 144'hf06ff6a9eed8036af55d0d8df4c6fdeef064;
mem[197] = 144'hf012fc02f9500c6ff79bfa5ff61cf86b078c;
mem[198] = 144'h0f7a079ff9bff9ecf1dc0e5903e505ce0f73;
mem[199] = 144'hf89ff187ff9bf47d0630087bf3f60272051c;
mem[200] = 144'h04580057f1a3ff8d0cce0ac4f6d4f9de0a18;
mem[201] = 144'h0539066ff02cff6d0cfff592ef540800f0f0;
mem[202] = 144'hf911f635f5010c130457f21406fef4a10e2b;
mem[203] = 144'hf56d0583f664080f0a5a0970f218fb5ef8c6;
mem[204] = 144'hfdfa0d31043dff74fb3a0073f3930c96f428;
mem[205] = 144'hff00fc7afc0f060a0340084ffb53f74b07fd;
mem[206] = 144'h069bf03afdd3ff6b0765fa1c0815faeef5a9;
mem[207] = 144'h0dfe026aff1bfb2df9f106d500ab0c690124;
mem[208] = 144'hfd760cf6f9e7f454f5a00d0f0738fd8bf153;
mem[209] = 144'hf28e0716f0d900cdf898f86b0693031cff24;
mem[210] = 144'hf148038a08780af40576f2f004c8f0cc0173;
mem[211] = 144'hf38bff19fe47f90df410f0780a9bfb10015d;
mem[212] = 144'hf545ea7bf659fe12f851edf809790322eff1;
mem[213] = 144'hf698f1b5efd0fadbf186fbf6f457f063f2bc;
mem[214] = 144'h0b0e06730b360474f6260ccdf9300136f701;
mem[215] = 144'hf567fe07f5d302050845f4a207ee024afaff;
mem[216] = 144'hfc99fb6bec7df7f80310fdb4ee04eec3f8bc;
mem[217] = 144'h02eaf08c0d61ef510139f4b5fff904c60c1c;
mem[218] = 144'h03cbffa9f9140d1a09cb0712fb53f85efbbb;
mem[219] = 144'h074efd82f304f808f663f35609d8fc9df844;
mem[220] = 144'h0cf0f582f170ee68ff19fc30fa39030d0a3a;
mem[221] = 144'h07eff3fa0cf6f396eff9ef9a02b2f2530327;
mem[222] = 144'h08faf84d041708a20b210b5901b3f0a5ffc3;
mem[223] = 144'h0289f3ebff1b08d7f30501270bb7f995f3a3;
mem[224] = 144'hf07601faee3b0cc103e90274f94ffbbeff5e;
mem[225] = 144'h090201c5ff7d0e9902d20bb60e40060efb55;
mem[226] = 144'hff14fdd808760e28000c0ef7f840fb52fd6e;
mem[227] = 144'h045a0a2df936f9280a51f473fc4afcbcf4c2;
mem[228] = 144'hf23effdc027602b5f01003edf8bdfecbfca6;
mem[229] = 144'h02e50b48f2faf2aa0b780002050a0731f94d;
mem[230] = 144'hf663faa8008afa850af00b18f31609d20477;
mem[231] = 144'hfe4d078dfd94020dff1300a7f8e7ff490570;
mem[232] = 144'hed45f5a1e61eea7ceb39f5f7f43eeb7cf2d6;
mem[233] = 144'h0493f9ef0b070b98fc8cedb70a240c1ffb72;
mem[234] = 144'hfab1f391efa8fa6ff53c07c5fe0bf56c0ac3;
mem[235] = 144'hf1240f5bf678f4f5f4a905a9f1ec09c3fd97;
mem[236] = 144'hf44ef31d099df9d2fb8004c2f886fb36fbb8;
mem[237] = 144'h0730f1e0f14a0deb06f6feb3ff95fd45fadc;
mem[238] = 144'hfa9f06bd0289ff98f7280b3d0a7efa4af027;
mem[239] = 144'hf803f9b008cc095bf3f80523f9c8eeeef0a3;
mem[240] = 144'hfa61fab3f1da05230713f92fff9ef798fc71;
mem[241] = 144'h0b190f80fde30ee1f8ebfbd9f95ff9b0fd7a;
mem[242] = 144'h0b1e0d53f75405cbf39f037cf7befb8f08ee;
mem[243] = 144'h0ce5fe99f01e06c1f90af234fb92018efcdd;
mem[244] = 144'h091bf318075e01aaf7be087af8fff6fd021e;
mem[245] = 144'hfbf708f5f99df8e204ac0c590510fc41f3f0;
mem[246] = 144'hfa4bf7deff14fac503b408600158f49a068f;
mem[247] = 144'h0731f3d8f162f6920060016d0259ef8cfbe3;
mem[248] = 144'h0c1907c9efa2f128fc79fb36fe13f873056f;
mem[249] = 144'hfffe0b51fdf3f7740e2df17d0b6e01700179;
mem[250] = 144'hf3ebf5f1f3ebf3120395fd850dadf7b6f0e0;
mem[251] = 144'h00870f990de1f8a0fd0ef55709d1f4410cea;
mem[252] = 144'hefc0048f0156f4be0610f81e00e307e40176;
mem[253] = 144'hfb40efb20b7204e3fa3d08b4f2080c360c33;
mem[254] = 144'hf5fb0c11f0fc043c0d82060cf5dd00cf0555;
mem[255] = 144'h089f090df20f0b1cfc6cf567fa76ffeb090a;
mem[256] = 144'hf44a01a3027a00df0a50f85cf835f3f60787;
mem[257] = 144'hfe61fc5cff7400930d57f44e0fd7099f05d6;
mem[258] = 144'hfcdbfcf8042401dffe970ca30216f894fc9d;
mem[259] = 144'hfaabfa1afc1b0565f0480652f0a907920c9f;
mem[260] = 144'hfcb4f2f80e9d0787f42404010246fa420335;
mem[261] = 144'h0592045a074cf443f394f2a20568f30efe80;
mem[262] = 144'h0ad1f741fe1b08d0072ff411fd81f4eb069e;
mem[263] = 144'hffb7fceef3c7fd34fbc5f585edb1fe26f60e;
mem[264] = 144'hf623ff41fcdc02070dc7f50af0ea017df7c9;
mem[265] = 144'hff9d03fffeb5fd9c0d30f0ad00eaf20eefa0;
mem[266] = 144'hf4f2f3cf0b250d9c01affe1ff395048df95e;
mem[267] = 144'hfbd1f24af863f3260ac9ff010e8606270275;
mem[268] = 144'h085909540489fec20c4f0b2efbbdf0f3048a;
mem[269] = 144'hf98b02a80a0afd1f084bfa400842fc500969;
mem[270] = 144'hff2307a207f7f9630ee20cdafefcf19d01bb;
mem[271] = 144'hf269fbc6ef36f56bfa4efac8f3140b700420;
mem[272] = 144'hfe6af994fe390bcbf09a0c7c0773fd66ff95;
mem[273] = 144'h035e0c31f53f0afdf02ef2a401bdf5b0f73e;
mem[274] = 144'hf7920bd1f83df4cc06fff636f1a30d3efb6c;
mem[275] = 144'hffb502c90023f8ddfbd9f23c08ca03c2fe99;
mem[276] = 144'hf193fe1e034d072308ca0f81fb060757f1f9;
mem[277] = 144'hfc5ef99b0d04fbf708eff5baf53706a2fefc;
mem[278] = 144'hf2200dc9fad2f741f475052206af0201077f;
mem[279] = 144'h0ba6fd2f0121ff62fe190d08fb100a51fd9a;
mem[280] = 144'hf8930fb8f0b50c5009e0faab0417fee3f449;
mem[281] = 144'hfa62022f0533fae0fe130e020cfd0303f04c;
mem[282] = 144'h066b0fd7fb0dfc27f520031bfb8af83afbb4;
mem[283] = 144'h080dffc9f4ddf3590a38f1bb02b908ad03c3;
mem[284] = 144'hf348f69b0017050005550a100d520df0faa9;
mem[285] = 144'h0639f3cb0b19064d0e2608a5fe980b9a001f;
mem[286] = 144'h09bbffd002440f4df6650bf00f29fe520f1d;
mem[287] = 144'h058b047d04710207f985f46f0865f2fa0d93;
mem[288] = 144'h0250f4a90b79ff95f5dbfbabf3a0fec1f9b8;
mem[289] = 144'hfb560c76fb410c6701e3079704faf7570eb9;
mem[290] = 144'h012f0572f1770ee50e900f9909b7037c0452;
mem[291] = 144'hf733042df3c50b31fbe0ffe3fac1f8dbf283;
mem[292] = 144'hf988fc7df070f8e0e9cd077e084fead9df58;
mem[293] = 144'hf32fef3ef5ec017bfa01fd9dfa83017f075a;
mem[294] = 144'h0972fe1ffc7ff1e00f7f02fe049b014cf2f0;
mem[295] = 144'h09d3f749fe51f9dceeff03c0f4e6fb5a08f8;
mem[296] = 144'h0617fae7f71fe052ef89f9d6f4f9e732f4ef;
mem[297] = 144'h0c720b9e0aa3f986f8f300ed054c0cb0f67a;
mem[298] = 144'h0e0206f70627f1e707e6f92df293ff87effd;
mem[299] = 144'hf8b40f4d04d900850fa00467f6440d5302b1;
mem[300] = 144'hff6904b7f07fee98fe0d066ffca00bcc0c1f;
mem[301] = 144'hfd11f09af8e80e0c07d3fcb0f63d097df68f;
mem[302] = 144'hfa06f61ff1a60f15f5ce0ae100cff4c8f365;
mem[303] = 144'h02f3fbeb09d6ff720ba608d803a4fe8bf71a;
mem[304] = 144'h095104c8f1f3eea7fe32f4c00793f938ef53;
mem[305] = 144'h0849fc400c010d9efbabfbdb0e2802aa0ebc;
mem[306] = 144'hfb9d0d8cfb0408f400e2f7b8f0aafb01fae8;
mem[307] = 144'h0865f066031ff20c0ae20827f5c608e904b5;
mem[308] = 144'h0ada0b13ead40622f8f1044cf618f7a1f6e0;
mem[309] = 144'hfa78f0c0f98b045af85af99a02b9f4e8fce6;
mem[310] = 144'h06b6082efc650dd90569fdbb0e1f0bb7f411;
mem[311] = 144'hf652f8a00465058eeb9509a0f60709250503;
mem[312] = 144'hed0ef9aafbd0f8c5ed84079ef2e501cceb7b;
mem[313] = 144'hf125f607fcf3f739fd52030f03690c000e0e;
mem[314] = 144'h0a43035bf729fa31fabb053c01010426f1cd;
mem[315] = 144'hf349022ffd39f6840569f7a5018c0d2af04b;
mem[316] = 144'hf0b40a630a980376088607bbfa38fe8006ae;
mem[317] = 144'h0e3b027c0c3bf6e6fec30b77fe9401dbff2a;
mem[318] = 144'hfa3ff9e3f715f5070b7e09a6fa8e06daf1c7;
mem[319] = 144'hf55ef40003a302a50e3a00cbf5540076f11b;
mem[320] = 144'hfd63048ef7e8fc16faf80dd709cc03e7f37a;
mem[321] = 144'h02d8071d077dfe47fb91fc08f7260ae9f863;
mem[322] = 144'h07fdfd36efeb0be50c8ff721f7dd010ff504;
mem[323] = 144'hfcd0f0910dcdf0f50c8df082055106b30d74;
mem[324] = 144'h0c2bf83eea3ceb5bfbf3e94dfb1e058cf474;
mem[325] = 144'h097f0214f02df18007d00c0ef39afcb407c4;
mem[326] = 144'hfb50fcca02bcf1cb0c840707014e02400219;
mem[327] = 144'h0b020679f17506f806e40969ef2cfad30a7b;
mem[328] = 144'hee06f882fa67fe37ea9dfdbafc4802060291;
mem[329] = 144'h0302078d0652ef4d01920737057803defa84;
mem[330] = 144'hfa23feb3033eeee80805f2d7007efb2cf254;
mem[331] = 144'hfc00fb190342f388f2cdf6c3faa6048bf6f4;
mem[332] = 144'hff430e11ffbff823ee92fc7d061df1fdfa6f;
mem[333] = 144'hf248fdf500abf14d046a08090e14019af89c;
mem[334] = 144'hf49ffa6eefd6f300088501c5f830064a03ca;
mem[335] = 144'h0091faabf502091dfe48fcefff3df96cf210;
mem[336] = 144'h010308fd00bf085afa8c04d0076ffc9fff09;
mem[337] = 144'h03850cfefcfb07dbf06bf99c0f4209a0fa17;
mem[338] = 144'h0879fd41f201052c0fa2fcddf90b017ff0c3;
mem[339] = 144'h0eb3f169f2300e25f77a0490f5c3f6a3fc9b;
mem[340] = 144'hfcefee6efe6802dbff0afdcf06d7087ef307;
mem[341] = 144'h062dfef90810f4a70bdc0b39f4200539047f;
mem[342] = 144'hfcec0633f260f198f7930e7bf210fef2ffd1;
mem[343] = 144'hfcabef9a0b76f79d01cdf4a807710a44f119;
mem[344] = 144'hfc1ff671eadef3a7f8bef137f80f0512f37b;
mem[345] = 144'h0a2cfaa8f3cbfe4e0c9d028507600a01f23e;
mem[346] = 144'h025200450b05f8220b91f368f8faedd50b56;
mem[347] = 144'h067cfb21f42d083bf50b00fbf4a70592effd;
mem[348] = 144'h0a9907def7d0f03b0bfe0257f9e40657f3e1;
mem[349] = 144'hf5d20ce40b6ef076069c03a80bb4fa00f167;
mem[350] = 144'h052ff571035cf982026308110ea50467f0b2;
mem[351] = 144'h07530e7e041e066a00e1f54d003c017ff09b;
mem[352] = 144'h0d9ffafef21c05d2f1e30f6efac8fdb8fc19;
mem[353] = 144'h0afa0cea0cff0e0605fdf96cf57502d80f73;
mem[354] = 144'hfb09ff96ffc4f918fee408fd05260f0cf728;
mem[355] = 144'h0395f1d5f92e02fa0205fda2f386ffd6f6ae;
mem[356] = 144'h0bb4f9b8f70105cffd8ef0e0fc28ff87eb39;
mem[357] = 144'h01d0fddcf4550cb7f7d60f7c0988fdb2eeb8;
mem[358] = 144'hf21c0553fc8900b103b8f1f9fdb3f962040e;
mem[359] = 144'h01f5fd28f0a9fcd8f398fd1ceb43021c0054;
mem[360] = 144'hef94ea8bf4d7f2ecf02004220aedf9a9e494;
mem[361] = 144'h056b0c5406530ccb0e32000b07c9fea90475;
mem[362] = 144'h0b92fc3deeaa09090138f7b8f961ffaa0716;
mem[363] = 144'h02fafde509890c5a0c6bf1cef5aff6a8f2dc;
mem[364] = 144'hf253f38e0616f770f3f0f18b00edf19f008b;
mem[365] = 144'h03d1fae9fbecfc56fab003b0fd740bc9efc9;
mem[366] = 144'h04390fc7066d06da0b490d4b0678f12b013b;
mem[367] = 144'hf6e30ce2f740fc7bf63c0d69f314f87e0406;
mem[368] = 144'h0cc4f7ef0cc702390858f63302af09530cbb;
mem[369] = 144'hfe9df287f2d409c501a7f8490e1cf00e0931;
mem[370] = 144'h0ef100bbf6b8076afba40ada0403086e0cda;
mem[371] = 144'hfb50f24600da0872fa41fc820e23f47b0be7;
mem[372] = 144'hff55f05ff48e064a058bfbcef79af580fc94;
mem[373] = 144'hf89a01b7ef9c06430b27f5e909f90c04f2fe;
mem[374] = 144'h0ab30d230c830f20fd78f8aff9d4fb500ce1;
mem[375] = 144'h03b6fc770de908faf549fde9f3330e9cf8eb;
mem[376] = 144'h04380aecfd41f7e9ff67f16508fcfd76fc75;
mem[377] = 144'h0d3bf7a300c4f8b40ed9feff0427f3e709db;
mem[378] = 144'h0a2d009c06baf6740655fbcd022cf60f0aa8;
mem[379] = 144'h0ce9fc9a08a4f41bf29afef50da9fd1305f1;
mem[380] = 144'hfaf90222f22dffdf07b5f924f6c9f381f646;
mem[381] = 144'hf6a4f084073801160c6cff55f547fa33f199;
mem[382] = 144'hfb850446fd820d180853fcf205120bdb00d4;
mem[383] = 144'h02c10600f669fd1d017805dc0f2bfee2f7d3;
mem[384] = 144'h016efb08041df006fcdc0a77ff000a14f1b3;
mem[385] = 144'h0c3ef10ef5b60dab0864fec40e9f0e360968;
mem[386] = 144'hfb62fefef0c3f8d6f2e4fd1a06cb06f10f6c;
mem[387] = 144'hf6ab0edcfe4bf440fed803360b5cf4020e26;
mem[388] = 144'h0d0cfe910084fb5df305f1f6fc8ef1bbf2d2;
mem[389] = 144'h024009580e41fd5cf1ab09c30b9cfb0cf8c9;
mem[390] = 144'hf96f0783ffbbf15afc2d021007460a35fb18;
mem[391] = 144'h0478f7caf4310677fb30f27a08250028f56e;
mem[392] = 144'hf0870b29f6940507fc95f7e3f084efc0f1e3;
mem[393] = 144'hfdfb0199f3d60c6cfd3cf7dd00d407f9f475;
mem[394] = 144'h0b5efa540f18f1230fc6f34909a003b6064d;
mem[395] = 144'hf2c70807f51507c1f335f146085ff33c018d;
mem[396] = 144'hfcf2fa17f759fe3cef81fa5b056bf462fda8;
mem[397] = 144'h01dbf93b00faf8aef0b6fc5df563fc4f08df;
mem[398] = 144'hfd38063d0f310ed8f315f2ddfd9ffea2feba;
mem[399] = 144'h041100a9007a0265f51209cb0676f32e01a0;
mem[400] = 144'h0ccdf9c10aaa04480526ffc6f2b20782fb7e;
mem[401] = 144'hffc902220dfcfdf909100f7cf59208d50384;
mem[402] = 144'hf5f20d630c4702ec0aebfce0f8b10a0dfe8f;
mem[403] = 144'hf254f1ed0cc7f89506600ef00b1a03acfb67;
mem[404] = 144'hf7500a69fa94fc6bf0110606f4de007dff94;
mem[405] = 144'hfb3a076d0a8cf07f01f60254f2aa04e2fd35;
mem[406] = 144'h0c8ff9be0cbbfe460cab089ef5d2ffe2fcf8;
mem[407] = 144'hf75f04cafe07f15300a709b2f8bfff9dfaa6;
mem[408] = 144'hfd9804f0e6f8f28dfbff0bb0071ddff3dff3;
mem[409] = 144'hf5e90868fe65015c08f20273fd42043d0ba6;
mem[410] = 144'hfe6ef597f5c9f790f831f596fc30f80b0474;
mem[411] = 144'hfebbf8b8f78cfe37fe910c1b080e08c80195;
mem[412] = 144'hef3e0abef3de08a1f398f320f24cfd55038f;
mem[413] = 144'h0e9efb2507200b1104beff54010202f4edf7;
mem[414] = 144'hfb47f34809b2fed3f29b0df30c2108e10083;
mem[415] = 144'hfc920476f1b7fe400e5efc2bf34bf0bbf622;
mem[416] = 144'hf1960ba6009df95aff8602cc0a6b0783fd92;
mem[417] = 144'h03dff00df2e10a17f792fc24f1affc5d08ab;
mem[418] = 144'hf22d097d03d4f6a8fd1008b10f86ee2af112;
mem[419] = 144'h0249fd190486ed0e02c2f261f353f1160670;
mem[420] = 144'hff9c09b60442ea11f70efccefd04ef41fa80;
mem[421] = 144'hf398f077051bf927099ef65802a0ed4dee9d;
mem[422] = 144'hf97b0b71f402086d0ab1f72ef47b013207f5;
mem[423] = 144'h00d6f351f1e9f166f24dfa720855f70ee51c;
mem[424] = 144'hf535fa4af754f357f50b0523fd06f36def29;
mem[425] = 144'hfc0d01c80070f329fe61f94dfd17f311fb74;
mem[426] = 144'h04e007eef786e9430426f7f50585f41b0974;
mem[427] = 144'hfbea0a87098f06a8f8140e51ffc5ff46ef9a;
mem[428] = 144'h032209a00bc6fac7eec80503fa57f2260e2f;
mem[429] = 144'hfc520827f05efb53f28f0e480b2c0838f4f3;
mem[430] = 144'hf3260104fb2cf7d2fd9c02b40403089602bd;
mem[431] = 144'h0498ef61fa26ffdff49af466f50205ddfe01;
mem[432] = 144'h09df081ef05c0507f19df16a05effff5f436;
mem[433] = 144'h01fdf657fc5e0f86f64c0e0ff8930bebfe49;
mem[434] = 144'hf9fef9b30f6800920839f7f8f99702370059;
mem[435] = 144'hf86f0e97079801c7f1f9f63af74cf657f30d;
mem[436] = 144'hf7d1f427fe520da6faa00f0903c60511fe61;
mem[437] = 144'hf097ff91f59c0315f37d093c01d3f0320344;
mem[438] = 144'hfcfcf93bf94d0aa40164ffd9f73f07d0f957;
mem[439] = 144'h00a1f0aeffeaf729f06b0c49ffe7f76df8b8;
mem[440] = 144'h0f20f5ae01bbf44003aff79bf2b6f3f2f14f;
mem[441] = 144'h0bc0f7c2fe4ef0280227f631ef9cfe4f077d;
mem[442] = 144'hf5d50cde0cc3fa7afc750c770d0df2b0044e;
mem[443] = 144'hfff608e60c3807fbf657f13cf508fde3045c;
mem[444] = 144'hfa8ef9bfefcef931fa37f35df0ef0a47f03a;
mem[445] = 144'h0909f397f1b60a6e00ecf205f5fcfc9cf445;
mem[446] = 144'hf9e604a0f171f1e209bcf7790128023f0fc3;
mem[447] = 144'h02d90edd08a6fba0000e0c98f9b604ac0329;
mem[448] = 144'hfa9df7dff84b07d9f98e01d4f7d4001f00d5;
mem[449] = 144'h0701f02ff8b6fb78fb7ef5400141052109fa;
mem[450] = 144'h0e6605f00e4f078701670bb4ff770ecc0fa3;
mem[451] = 144'h028bff28034f0c470c420b8309b0093cf5a1;
mem[452] = 144'h099cf56608aef50b07210a45f5bc076df011;
mem[453] = 144'h0c4bf03ef35107430b39fc9909f2008d0381;
mem[454] = 144'h0b0d0c4009eef5860974f6b5f55003100140;
mem[455] = 144'hfa200325fa610699eeedf3910ae9f093efbb;
mem[456] = 144'h043ef39f0422ef5cf0c2fb1604f80997f031;
mem[457] = 144'h05980115f7a304acfca5ee7cf7e008bbfcdf;
mem[458] = 144'hf3a0f92cfd90fa2e04a30759f1e3f09ef4fa;
mem[459] = 144'h0e6901c2fc6507aaf7b40bb403c001e80316;
mem[460] = 144'hf80c08f104ee048e0a070bd20d130aac09a8;
mem[461] = 144'hfd64fa30f8810ec00395f309ef31f38cf62d;
mem[462] = 144'hf262f7d30bbd015ff6eefaf206ba01a00bf3;
mem[463] = 144'hf0e80851fd7c0083021b03be078601d4f08a;
mem[464] = 144'hf749027ff2ee09890ee104450ee703980b48;
mem[465] = 144'h01750938f23bf56206f60d9108c4f78df3b8;
mem[466] = 144'h04060aaffeeb07c8ff3b05d4f3dc00d7085f;
mem[467] = 144'hf102f603f023fd8306b2f1dd093601f8f1c6;
mem[468] = 144'h006b0bfc08460094f28fffbd0b6906020650;
mem[469] = 144'h0a1709d7f716f54d02bff39006d50a2efa64;
mem[470] = 144'hff180f5208e7fcf7f2e90f11fc780f680a35;
mem[471] = 144'h02c7ee390329fac5f669f68e0aa70a33ef3f;
mem[472] = 144'hf4d3ef7405a8f23ffc73f4b8fccdf89bf5b5;
mem[473] = 144'hf923fb10ff28efc0fcb40c6dfa89facffe5a;
mem[474] = 144'h0f12fa5ff0abf1f50736ff5ef335f82d0b28;
mem[475] = 144'h00140be90272088405cb041d08a202d10258;
mem[476] = 144'hf905011cfb48f14a08430b60fd82055904e1;
mem[477] = 144'h077cf53ffe96f32bf14b0827fbf40ec8f9ed;
mem[478] = 144'hf0e00a2803670200048900480a5ff033f500;
mem[479] = 144'h064e083dfe31f2430a17f7ccff49f79b0bb3;
mem[480] = 144'h0a4d08790411f0da0db7ffecf5b5f2e3f638;
mem[481] = 144'h0915f604f6140a33f3eb08180342f5390036;
mem[482] = 144'hf6a7f9d60f99fce8f8870f460cb2f1fe0ee9;
mem[483] = 144'h0caf0fe80470fb10fdf2f292f8a30558f026;
mem[484] = 144'hfafc082f003cf046fce4f16806d90bc20dfe;
mem[485] = 144'h0b5d0b9a034109dcf10601c7f095024af861;
mem[486] = 144'h000efec30d700cb8fae4f96befd005cdf299;
mem[487] = 144'h05e5ef21f303f883024d0340016205fff8fb;
mem[488] = 144'hf9cdf23c0016fc13fcd90686fee409ac0104;
mem[489] = 144'hf18d0f550180f6f5f32f031c0bf10e820dc5;
mem[490] = 144'hf1dd007cf8a70d61f0980337038d03af05f6;
mem[491] = 144'h0658f3bdfa0807f804bb08db06a8f2c4080d;
mem[492] = 144'hf65d0576fd2f0a80feba0e7ef53a08ac08d6;
mem[493] = 144'hf38f0a08f1470d53f49a09eff0d208740ea4;
mem[494] = 144'hf8030081f208fefef9c208e6f8310f84fd47;
mem[495] = 144'h09e20de1018efb31fc22076bf72bff230313;
mem[496] = 144'hfb230b11f1ec08e5fc14f1e8f999f7dcf4f3;
mem[497] = 144'hfe480e75fd5a02c8fdc00b69fa1d0b8e06e7;
mem[498] = 144'hfaa7f5030b49f525f454f5eff79d020f0dbf;
mem[499] = 144'hf59b0f09fa310068f58102bff9f40edd0086;
mem[500] = 144'hf838036000b00822088005ecfa3cf7bc0b67;
mem[501] = 144'h08120c840e20f71bf10bf4160b4f0e770c54;
mem[502] = 144'h05cf0b3ff6c6fc99014a05f2049a030802c9;
mem[503] = 144'hf53ffcd400b2fd94fd96fc05f990f20b0a1e;
mem[504] = 144'hfb6d06befabcff95f68e0b95f5a6f0c600f2;
mem[505] = 144'h0424068f0c6ff588fc7608d70e91f55af510;
mem[506] = 144'h0fc1f6f0fec602b702d8f079f3ebf88df912;
mem[507] = 144'h0a290b6a075e076afc5dff000d870f9cf443;
mem[508] = 144'hfda403bef14bfa62fc7001420bbaf597ff3b;
mem[509] = 144'hfff00ba8f39a0b1100ecf677f831012cfccb;
mem[510] = 144'hfb72f08df755f9d601d0f4caf5b1fb3f0501;
mem[511] = 144'hf39a0dd70bc2041e0834f3e7f453f788024b;
mem[512] = 144'hf54b0cd5058e021b0393007afcf8036af1e8;
mem[513] = 144'h0d2c088ff9460eacf068033dfdcafa3ff7b5;
mem[514] = 144'hfaf4f268f9e2f0a6f277f6eaf20ef749f77c;
mem[515] = 144'h07110582f323f2d0fd18f105fbd5092cf783;
mem[516] = 144'hf526096b0478f91d0b35f1e308a109540957;
mem[517] = 144'h02c60323fdc80c3bf319f63bfe18fa48fbb3;
mem[518] = 144'hf8d8faa2fb5102a8fe24fbbe016a0805092b;
mem[519] = 144'h0871eff8f07ffee208ddedb709ca037cee51;
mem[520] = 144'h08bcf4d9f93cf4e4f90bfa1d069407f7f9fe;
mem[521] = 144'h0bf9f059f3f0fd91fbe2fc68f728fc300653;
mem[522] = 144'hf6a20e00fc27069dfdd9f6ed054a0b2206a5;
mem[523] = 144'hf9c30d3c00d0fc5a0f410f0c042f0476fe78;
mem[524] = 144'hf25f0c080502ef9cfc55038e01d001110856;
mem[525] = 144'hfa0d0cdd0d84f2a505e00f2d035dfb0a0173;
mem[526] = 144'h0c62f5a5049df4ba0c2e016409ff0841002e;
mem[527] = 144'hfadb0abd023dffbd06d507b00b45f2c7f551;
mem[528] = 144'hf0d901abfc9af0b60031f15df695f615020b;
mem[529] = 144'hf2b209c50631ff61f1e4f3240ab0f96f000f;
mem[530] = 144'h0c2505dd0d47f1c90a6cfa03fa83fc90f22a;
mem[531] = 144'hf3b3f194f193071eef38f268fc370615efeb;
mem[532] = 144'h01b4feb6fc6af325ef23f6dff86ae773e973;
mem[533] = 144'hf4e302b1f52c0acd0660fcb0fc0cf6f50297;
mem[534] = 144'h0a12f24005d2fa39f305fc320c5800c8f152;
mem[535] = 144'hf35fee9bf7affe0ffd1b066f0660086a08c1;
mem[536] = 144'hf39cfd850032efa4f2f6f228ff13fe31ea11;
mem[537] = 144'h05ddfbecf81e0176f4f6fc5b0a9d08b3006b;
mem[538] = 144'h0aa5f13df5e9044ffed5fb8feec507650575;
mem[539] = 144'h060ef73606030fd7f66e07a9fea2faecf1cf;
mem[540] = 144'h004af53707edfb900a9d0e1bf0c2f3bf0359;
mem[541] = 144'hf26d06b402fbefb90ee905f50e40000eeff5;
mem[542] = 144'h051efa9cfb95fec7fc12fc480c39f6bcf0ae;
mem[543] = 144'hf17fefc6fb4201f80e9d0233f4290ae3ef41;
mem[544] = 144'h0e86f0caf6dbf6760a590ae2f60a067beed9;
mem[545] = 144'h0feefd67f70cf77e063bfe4103f5fc61faf5;
mem[546] = 144'hffc1ffb4f2d40d7bfac708100eb7f288fc95;
mem[547] = 144'hff25f5ea0b6bfaf2005ffba5f12007aa051e;
mem[548] = 144'h09550a84f1c1f06b070701b00464fc01f5e1;
mem[549] = 144'hf6c2fa47ee34fe5fffd0fec9fe6004e0f89d;
mem[550] = 144'h0fb60f2d0d1ef8990382fc0d00970881f7de;
mem[551] = 144'hf112ff4d00a6f291066c012ff4a30407f6fb;
mem[552] = 144'h011ff6a8014d04a8fd36f4c6f790f23df630;
mem[553] = 144'h0a21058f07930012f92609dbf973f64df520;
mem[554] = 144'hf9ac003cfe16efb6f86f063afe2cfcb4f6b7;
mem[555] = 144'h006e0e3cfe16f09f04630498f4df076e0718;
mem[556] = 144'h0081f0e9fea704fafc42ffe70b55041f0068;
mem[557] = 144'hfe2200f8013ff83ef102ef0df506f253062b;
mem[558] = 144'h0637f39801120aae08d1f527f4d5fd640c46;
mem[559] = 144'hf8a8f10303d6039404970c7dfb140892ff32;
mem[560] = 144'h05a8f612fd7ef1650d5d02a6065ff6a7f5c0;
mem[561] = 144'h0741f9760e4705430948049ff897074208e1;
mem[562] = 144'h01ccfd03f137021f04edfbc4f5d5f088f2da;
mem[563] = 144'h07a5f12bf789f3f4016afffc0d66f709ff34;
mem[564] = 144'h0a0d08a2f283f212e69c01fef780fcf4046e;
mem[565] = 144'heefd05c8ee90f697f211f4e0fb35f22e071a;
mem[566] = 144'h07f5f895fdcdfb6d049501a0f49a0d03f178;
mem[567] = 144'hed1af70bfc1b07c1fed200870852f19af840;
mem[568] = 144'hfbe2ff23e948eaa0fb39077ff455f7f709b1;
mem[569] = 144'h03f5f093fe36f63cfa7403a4f9b7f0fc0786;
mem[570] = 144'hf8da0879ec76031c05920123fc14006ef470;
mem[571] = 144'hff5df1dafc2c08dafed00ed9fdb0efe807bc;
mem[572] = 144'hffba0c72f48301c10d80fd35f1280eefff04;
mem[573] = 144'hf7a8fc63f4fcfb820decefe00e9c07e0f39c;
mem[574] = 144'hfaf504dc075f05a30d4d0d620bde008f032c;
mem[575] = 144'hf2da0e61f3da0774052901da0874fac00175;
mem[576] = 144'h0b730b180579010cf2320614f5b4f0b30edc;
mem[577] = 144'h01d2059df97e0d030cf5f1be0072f51b0524;
mem[578] = 144'h092a08dfefb60435f3570357f91b09740809;
mem[579] = 144'h0108ffedff21fb8cf169f67108f3fc980b33;
mem[580] = 144'h0a95ef56ffe50471f6f602f606c50aa0fae9;
mem[581] = 144'hfa24f7260a7af531f224f35dfb6f0e86f203;
mem[582] = 144'h0da70334031703e90259fa6ff58c0819f7dd;
mem[583] = 144'hff80f21108a1f85af90eee260492f03bf3ea;
mem[584] = 144'hffb9083806190462f49efadf05f1f38605f3;
mem[585] = 144'hf23ff84df623f8990cb9f06b0b9808ecfe2c;
mem[586] = 144'hf950fb3ff96b0dfcf2790e310c790380f7e6;
mem[587] = 144'h063002060bcd0c61fdeb01bc0997f153f858;
mem[588] = 144'h00abf30d0aa5f42f05e5f0220c93f04af32b;
mem[589] = 144'hf0ce02880209fef208150c060593fa0104bb;
mem[590] = 144'h0878f80c01d0032ffb2bf522f8b3f6e4fc63;
mem[591] = 144'h0eef0d43f1db01170742fbf10695feb4fed3;
mem[592] = 144'h0e0afce2098d01190c0804b00096f9100838;
mem[593] = 144'hf48b0b44f4bb03790ce7f0840c5505d70f36;
mem[594] = 144'hfb2ff6b7f9a1f01902cbfc450001f809fb23;
mem[595] = 144'h04510e1bfbcdf84ffbecfbc404a8f82a012c;
mem[596] = 144'hf746efc70ac809c0fc12f17d0711033d0e7d;
mem[597] = 144'h075bf309f334f18af84c0517f5ecf7abfa39;
mem[598] = 144'h06a50d1605b1fdddfdd7f7f20f7cf81cf93b;
mem[599] = 144'hfab1fe8d014c0b7df504f5eefa68f54b0410;
mem[600] = 144'hfaf0024d02b4fae6f93fff1703b9f2ac07c3;
mem[601] = 144'hf8e6fd550888f232041f047c0c80041bf7c0;
mem[602] = 144'h067df97b0eb8f90002ce0e62000ef778068a;
mem[603] = 144'hffddfd8c04a6f76ffa2a05dd0c08f7fb022d;
mem[604] = 144'h01c3081a0b2a0a990b54f1260049f99aff76;
mem[605] = 144'hf5a6fa8ff21c0709029f0f10f9e2fe9100a2;
mem[606] = 144'hf60dff230d5d0699013dfcaa0374faf1fda9;
mem[607] = 144'hfb8c05960468f28af78006770330f6bf03f1;
mem[608] = 144'h05c40520fa10f23001ff03f3f97a01bcf7c3;
mem[609] = 144'h0acd0be501c6fa510425f945f59304950dfa;
mem[610] = 144'hf70af9c6fbcdf6e0f3ac019d0428fff8fe5f;
mem[611] = 144'h0ea3027bf86cf99200280d3c0f30f6dd0ef0;
mem[612] = 144'h00430631f491fcc2fe0cf9780697fe92f89b;
mem[613] = 144'hf8fe0b410632f509f3230fabf360f4a8ffed;
mem[614] = 144'h049af857096f053105b20bb109560e52ff50;
mem[615] = 144'h0b70fc280f3f01c00651024f095b04d9f41f;
mem[616] = 144'hffd90b850c440c38fe49f709fc2bf906f537;
mem[617] = 144'h01b00bc30b5f0cebf1b50f920cfd0e3a0f7e;
mem[618] = 144'h0535f8c9fb2bf246fec60598057bffc40aeb;
mem[619] = 144'h04a604abffd7f0e505f50ead0d170fbd0524;
mem[620] = 144'h01bbfeef055708b1f4e50705fd5ffe47f9a9;
mem[621] = 144'h05bcfe43f8c402370395f907f416044d08f4;
mem[622] = 144'hf29c0f68fcc402cc020ff4c4005701af0516;
mem[623] = 144'hfbd90895fd65f7fd0fb0fe140b7f00260e3d;
mem[624] = 144'h0d5308b9f97e0e92f5610e68fec90ed80563;
mem[625] = 144'h072e0ca40930ff7ff4050dae0a3c0a390252;
mem[626] = 144'h0a4a0745f378f21ff7f2fc54fc890064f5e0;
mem[627] = 144'hf7bffdcef7a2efa90ad0fae1f3fbf8b80770;
mem[628] = 144'h053d04150b15f704fa780b99f695f38cfad8;
mem[629] = 144'hef550ed003ec034c0be70449060606dff329;
mem[630] = 144'h0d6efad80b32fed7f5e4f243fce50b6206a0;
mem[631] = 144'hfdf208460a6ffb5df9930aaef884fba5f899;
mem[632] = 144'h0020031502f2efd906e705e00d3e0ae2efc3;
mem[633] = 144'hf57f08f9efa4fbf0ef46f34bf434f5630603;
mem[634] = 144'h06bafb53fea6015afe84008df67f0440f2e7;
mem[635] = 144'h0ad4094c0a5c0ddbf7d9fa270c3a06fef3a8;
mem[636] = 144'h0df5f789f2370147f8ecff82fbd3046cfd69;
mem[637] = 144'h00a6f9f5f88a03f8f57f058e06e3fc17fd48;
mem[638] = 144'hf1610b08f3f9fd50f796074602a3043ffa89;
mem[639] = 144'h06e60076fc58061c0dcb09390a5d09fcef35;
mem[640] = 144'hf835f7d2fab5f7e4f70df5a90d9a05dff45f;
mem[641] = 144'hfd590ae7fe09fcdff1da0068f5cafc16f27f;
mem[642] = 144'hf266fe6806adf52afd40054b05adf07f078c;
mem[643] = 144'h041e030d0622f73a07b2013e006405740de4;
mem[644] = 144'hf2dcfe82f7080570f1460750f56ef88b070e;
mem[645] = 144'hf0980443f61f08050b50f6d6f058f4d90e9a;
mem[646] = 144'h083a086cfe0dfc2d0cd30b8df70f0299fc84;
mem[647] = 144'hf9c5f89f036cfe840081f5c2ff1dfe39f9a9;
mem[648] = 144'h05bcf06af85d0c7b04b6098b0f050a5df567;
mem[649] = 144'h009e0211fcb40c5b0d6203f4f3ed02dbf995;
mem[650] = 144'hf3400881006f0e600c17f56700daf0090665;
mem[651] = 144'h04d20a720828fe2ff401088d0562efd80885;
mem[652] = 144'h07f40479f9c60aa60a4201200d020aab0cee;
mem[653] = 144'h0a670e51f326fb21fc95fae90ee0f3050785;
mem[654] = 144'hf08003c8f3df00d6ffbb0fa20beafdfcf9f8;
mem[655] = 144'hff96081f070e060401810cd0ff0cf17ef3ed;
mem[656] = 144'h0c50013e0386f8a3053afebaf67804d90131;
mem[657] = 144'hf8b5ff3d0f9df26608870bbcf2fcf302fc9e;
mem[658] = 144'hf283fc090deaf21e0620f078f3a70ab6f578;
mem[659] = 144'h07d3f664f14cfe1d0754f4e20022fc5206a2;
mem[660] = 144'h00d0fc2cfa750035f3d4fa17fed902e0fa23;
mem[661] = 144'h054fef52f9d9fc95f42707f90ed607a8f9e4;
mem[662] = 144'hf4fc006b06effbef0f8c0aaafb9bf3a20028;
mem[663] = 144'hf717f73cf22afed5003ef216ec8bf33a06c4;
mem[664] = 144'h0c41fe0cf958fb29e8b4fada011bed28f31d;
mem[665] = 144'hf32506b7efc603080bc3fc430935f1250607;
mem[666] = 144'h058ef67809100c9d0475f05efec2fcf5f103;
mem[667] = 144'hfeef09820f8ef362f53c0454068afdd5f023;
mem[668] = 144'h0427fca505e40995f84bee9008b8f8200d11;
mem[669] = 144'hf8ac0ef1f4f1077bf3adff1a07d305eef2ec;
mem[670] = 144'hf058fa84036405ffffd5f082fe00f598f136;
mem[671] = 144'hf6240ae8fb7df6480cd40796fda00b1b0dd7;
mem[672] = 144'h0d6af7060ae7f96302f80af4effe01ab0b18;
mem[673] = 144'hfa0cff82fdc202b807a3fc17f0f90b64f522;
mem[674] = 144'hf9e1f7d8fa0cf3e10bcf0a05f22cfe7f0803;
mem[675] = 144'h0b47056e08dff4130aaefab5f4130164f749;
mem[676] = 144'hf95bf1d7f1df06210e5403b706880767017b;
mem[677] = 144'hf82f0969084af7a4f363fb8df1d1078e0e14;
mem[678] = 144'h0b03fb2708b10e8b0e14fee6fd8e077af394;
mem[679] = 144'hfe31fb23fb780135053df9a30ca2020df03e;
mem[680] = 144'h0697077808aaf89bf25af7abfe6af887f321;
mem[681] = 144'h04b402550dee0e22f0a1f928fc09081e0328;
mem[682] = 144'hf24f0c1afed0f1b3f154f11f01820982064d;
mem[683] = 144'hf849f175036ffaa5f091f0b207cafb6b09be;
mem[684] = 144'hfafcf97f03d7081909bf02d308e302b80256;
mem[685] = 144'h0efbfb63fc6df4fcf7ae05fafc82f71003b0;
mem[686] = 144'hfbe2fe98fee1f61b03600ceafb4efbf3fa47;
mem[687] = 144'hf1b6070bf9b2f4280ae603a705d007adf4f8;
mem[688] = 144'hf99af034085ff15802c2ffe70d0201110ccb;
mem[689] = 144'h029df217f9bc0c2004070c4df05306d20fdb;
mem[690] = 144'h0b600298093ff24c0a17fb32f1730f5bf7b8;
mem[691] = 144'h0577fa5df958fc05f7940b3d049cf66bf2ca;
mem[692] = 144'hfc3109cd0038fc4c09bd0850f008f092f25a;
mem[693] = 144'hf3260d5508b703e2076f0650fc8af2c40460;
mem[694] = 144'h0f67fb68fefdf533fa4008b0f25602bf051d;
mem[695] = 144'hf174f351fd520703fe05fd15feaa003e0dd6;
mem[696] = 144'h0676f79bef9af703051ff759f3800bd40973;
mem[697] = 144'h09b7faf5fa360a38fe460fc50f20079b0a92;
mem[698] = 144'h0c81f81c0e48fb1004700c52f476f97bf136;
mem[699] = 144'h0949f6eef474085bf413f2edf8250159030f;
mem[700] = 144'hf855f382fb46f7320c700da7f821fa23fad8;
mem[701] = 144'h0129f6d0fb3b0cc9f712fac20c520e20f995;
mem[702] = 144'h08ccfa6f01f205fafa3ffaf8f8cdfcdef89e;
mem[703] = 144'h008c0d56025c04e2f1def4d5083ef6c308f2;
mem[704] = 144'hf25908880c0400b00ef9086505c20c05faff;
mem[705] = 144'h060ffe9ff7e201b00750011b0ef5026600a7;
mem[706] = 144'hff2d09dd055af897f77006e501b90236039c;
mem[707] = 144'h0f00044a0ad1fe6cfab30ecefd08037a059b;
mem[708] = 144'h0115fbfaf25aefac006ff797f61c0b16f1f7;
mem[709] = 144'hfbfbf286089c0a34f7800477fa660f3bfe4c;
mem[710] = 144'hff9408aa03dfff4bf27f085409d8082dfd80;
mem[711] = 144'h01a4ff530b93fb8fefca01cd0c0d0275fc1b;
mem[712] = 144'h03a2fcc401b2fde904a0f7ec0ea300840603;
mem[713] = 144'hf3f4f0fc04ecfa1afe54ff4f0a12fae80b3e;
mem[714] = 144'h063402670de2ff24093bf76f0c3ff28d0c8a;
mem[715] = 144'hf476f55904e8fc32f6eb08edffbbf1690f65;
mem[716] = 144'h0e64f40dffa70431f3fa04820685f4a20938;
mem[717] = 144'hf1520340f9bff72bfcdcfd8d078af8830dc5;
mem[718] = 144'hfad8f8c802690974fe4e0b8cf5faf8830290;
mem[719] = 144'h058cf1a2ffbf07940159f5f7f0e9080c0af3;
mem[720] = 144'h088ef0b10bc8f8290293f5c1007afc8dff7f;
mem[721] = 144'h0ba4030d0eb8f985f66f0c8a0c6a07b50c53;
mem[722] = 144'hfa60f19df381f148fb150eaf0c810bf9fb10;
mem[723] = 144'hf017fb5fff7900b30ec801060620090c09aa;
mem[724] = 144'hfda50d16fb470e0d0925f69907890cbaf60b;
mem[725] = 144'h040a0d6efffaf63df215f0bd04b5055bf7e3;
mem[726] = 144'h0dd8f35805f50ee6f067f584f2b8f1e00b58;
mem[727] = 144'hf1fef312f3910c0cf601f1f70448fde20828;
mem[728] = 144'hfe1d0d9e0a06f21504af038ffebff608f2cd;
mem[729] = 144'h055c084e0077f41603980902fc03f4fb072a;
mem[730] = 144'hfdf6f2a7061c0c81f295f18bf3e9060ff793;
mem[731] = 144'h086bfaa4074702e80473f0eb0e860e61f6c4;
mem[732] = 144'h076ff45f073cf1a0062a0582fbd609a5fff2;
mem[733] = 144'hf6050ce6f0370a0100850555fc680dd0061f;
mem[734] = 144'h0722ffcff3b3f077018e0eb60ccb076ff7ab;
mem[735] = 144'h01b10d8ff4c90018fc83fe81f51a0f82f5fe;
mem[736] = 144'hf2b7fc7ff541fce2f32d061f00aafe8e05bc;
mem[737] = 144'hf6bff371f6fc0c8a095af344f1910812049c;
mem[738] = 144'hfeb5f4a2071f07cf0ebd003c02b4f7a80719;
mem[739] = 144'hf28ff4d7f746014cf4540c5f0632f1c5f472;
mem[740] = 144'hf7570a6a04fdfe84fe36f8f20fa1050e0bfb;
mem[741] = 144'hfa860beaf7da08e6fafcf925ff5bf8bbf551;
mem[742] = 144'h00f4f24ef5100d7c06b80ebf0c7cfcee0e69;
mem[743] = 144'hf4b203c40e990dbaf7370d51fd72f9ecfd01;
mem[744] = 144'hfd36fab8f4160cd4fe5bf28b04e40a82f1f2;
mem[745] = 144'h056cfb730ef90823f577fae1f79e0b1ffc47;
mem[746] = 144'h04e90031f608fecc0e3df4d3f50a08280157;
mem[747] = 144'h08800624fe6c0004fe06f3b3fc6f046dfdcc;
mem[748] = 144'hf4a305c0002c0c58f48dff4f0396f6c7f721;
mem[749] = 144'h068b0b22090303510ca902110a5b0217fcfc;
mem[750] = 144'hf803f8adfd00ff1f015601eb050df9c3f01e;
mem[751] = 144'hfc520c24f863f2bc053f071f05390490fda8;
mem[752] = 144'h0752f8140b350e52f5540d42f34bf6a90688;
mem[753] = 144'h0037fb00fca8096a0f2ff6c9057201c3feeb;
mem[754] = 144'h0592ffb90c3e0e3cf9a405510102f3c3f3c0;
mem[755] = 144'h022af2b4f70efaa2f35007fdf9a80fa4fa09;
mem[756] = 144'hf0e502eaf0cc0c4402ad08e1f64af1400581;
mem[757] = 144'h042ff7c20330013afd890cfaf0bff89f02d8;
mem[758] = 144'h06650eaaf8a4f06d0ccd0c2d0c240c7af7d2;
mem[759] = 144'h002d0e99f71e0270007bf5f3f2e40c90f602;
mem[760] = 144'hff8cf1f1fa9ffcb10e1afa08f13efa2af07c;
mem[761] = 144'hfd80f340f7c80e040a5708f2fe54f100f229;
mem[762] = 144'h0e550eb2f05d0db80918fb79fd54f2200999;
mem[763] = 144'hf2b4fda5f82e0955f85af232f998fccafecf;
mem[764] = 144'hf791042609e2f951f34ef0d0fab8f32c0828;
mem[765] = 144'h05c7f29d02f9fc60fa67f37307930a40fa3f;
mem[766] = 144'h029e0b49fdac0fa7f806f443fdf6ff5cf400;
mem[767] = 144'h00a4fd0ef773fc530f3009a5fa9cfc65f818;
mem[768] = 144'hfe54f66f0e710d1df342f5330fe60824fea1;
mem[769] = 144'hfd9af871f71d08bdfd5b06690f4009a0f301;
mem[770] = 144'h02580c6befcef713f4effdbe0499f4d3f5c9;
mem[771] = 144'hfacc0795f9aff6560caff4470a870373fed7;
mem[772] = 144'hf0cbf26e02fc099a0e2bfcc9f76fff5302ac;
mem[773] = 144'h0461fc0100e5ffa9ffa0049af0c1ff91f48f;
mem[774] = 144'h05e40d000002f091042a0339f3640ba707d8;
mem[775] = 144'hfdfc034e05b4f97af6d90d350d2df9abf10a;
mem[776] = 144'hfd960726f418fbe402a4f81003850b76fe39;
mem[777] = 144'hf83a02cc0809f0050214f4e2fbbffed5f4e6;
mem[778] = 144'h0892f5b30c8df063f72d0791ffe70e4f0cb8;
mem[779] = 144'hf666033c0bfe06260b84fbec095affabfc15;
mem[780] = 144'h00140e25027bffd90de2f17fffe609440da6;
mem[781] = 144'h0907f6ccfd7bfcd8fd2a08cd049c0447f753;
mem[782] = 144'h0da7f922f43dfe650b0c0264f157f364ffe6;
mem[783] = 144'hf04d0bd5ff250521f6d3f0b6fd82fc2afcf5;
mem[784] = 144'h04d3051a0890f3b3f489fdadfb73016afb88;
mem[785] = 144'hf7a60281f895031bf7c6fb87f70a05690ede;
mem[786] = 144'h0af6fa00f326031d07ca0b2ffd0af1dff61b;
mem[787] = 144'h036c0ab90f9ef486f370efe008940ef8061f;
mem[788] = 144'hf8acf7670c360a970620f2e9fa9a0595f0d7;
mem[789] = 144'h0cd2f2d6fac5011b0692f944fc7501dbfc36;
mem[790] = 144'h0ebafbc0f671fdd8f8a0f0a0f2250de90ed6;
mem[791] = 144'hfae007460924efb80350f96ff712ff2f0b15;
mem[792] = 144'h0359f55bff6df020ef93fead064100c4f28c;
mem[793] = 144'hf386f6da043d0d01031cf8b20b81f5ea0efe;
mem[794] = 144'h0c1b0b36ff9bf175fbc30a6b0abd037b0b8e;
mem[795] = 144'hf9c60ea30611079ff22cf3e6f600028efc64;
mem[796] = 144'hf47e02adf000026defa907a60ab3f01108cb;
mem[797] = 144'hf07ff2b904820eff0671fdd7f7fbf5fef695;
mem[798] = 144'h018df666f1e00497ff83ff87f54cf58106b0;
mem[799] = 144'hff9f08b803650262f8baf87404050cc20717;
mem[800] = 144'hf5680b6b098e02120517f13403defa1af82c;
mem[801] = 144'h083dfdd1fd3b01acff46f007f2a500b9029b;
mem[802] = 144'hf1cbf6cdfaf4fda3f8d904edf815f5fefb5d;
mem[803] = 144'hf3c7fae4f51c0115072908c50edf0a4801bb;
mem[804] = 144'h0576e8f7f32cf2def643f4eaf219e7fff68f;
mem[805] = 144'h05900a01f1adf87c0bc40192fd34f44102f1;
mem[806] = 144'h06cbf2cdfe45f194f609f5c9fd5ef96e054c;
mem[807] = 144'hfef3f8aef512f6fbff510974f486f020f7ad;
mem[808] = 144'h07530043fa04f2f9e170e9a4fa21f084fb7a;
mem[809] = 144'hfcfa0e39f0110acdf1a00097f5f5f6d6f698;
mem[810] = 144'hf9affcbdf426f4dd0a8805080d5efd960254;
mem[811] = 144'h0147fe23f91a0eb20105f156f5ac06acf824;
mem[812] = 144'h0acd0791f6a2f47bf5fcf0a100a0070d0727;
mem[813] = 144'hfde3ff630bbbf8b80aaff52cf9e1f614ff0f;
mem[814] = 144'h0b0801430435097809b9f0b103f0060e0741;
mem[815] = 144'h0d460c85fcd406cf0ed6fec4eed00142048d;
mem[816] = 144'h00f9efd2f187fb36045df734fc880616f1ed;
mem[817] = 144'h094dfd1f0fadf94d053bfc39fb7105cff4ba;
mem[818] = 144'hf83af1b80cfef579fa7c0021036b0b76fce3;
mem[819] = 144'h0297f3e20ab5fa0d069d0023032bf02befda;
mem[820] = 144'hfa32f2f908cff8a501ac0c8afa5ef6b1f74c;
mem[821] = 144'hf2a2f40cff12fbf80572fb180d9801b80531;
mem[822] = 144'h079cfb9a09950b4c0f4df96c0c0bf27102a3;
mem[823] = 144'h049df16c0bec051104f8f06dff5c0b8e09ce;
mem[824] = 144'h0372fdadecd7fe29f01f080006ecf0d00271;
mem[825] = 144'hf7830b83ef19f915fc1af49ff5d5f0900d48;
mem[826] = 144'hf958fd8af5a7f36407dc06ac07faf02ef9c2;
mem[827] = 144'h0d14f8190610025d0c9802e1f644059ffdf2;
mem[828] = 144'h0600fb6ff16908cbf3fd032d0c4cfd670af6;
mem[829] = 144'h09f5f0d5f7cbefe0f5ed01be005cf4c30422;
mem[830] = 144'h0c68f66209290565fc11fed306e8f0ac08d1;
mem[831] = 144'hf8a9ff9c0acef946f888fa22ff180c82efa3;
mem[832] = 144'h0441078c044606cbfbdf0551f016f2f8fded;
mem[833] = 144'hfc50f19b0cf1014b0b20fa2c07750e84fcaf;
mem[834] = 144'h05e0f1bc0fe5f638f00afbca04200899f731;
mem[835] = 144'h0bbaf2380aa50480f389f70efb77fda00e3d;
mem[836] = 144'h07a80a7606590268f286015b00d7f7cdf4ff;
mem[837] = 144'h054eff3ef4460c6d0902f51cf84cfceafd69;
mem[838] = 144'hf8ec05e805600a33fd0801460241ff72fed2;
mem[839] = 144'h017dfcacf9bb0069f576f4e50a6909beff7f;
mem[840] = 144'h037e047f0cbef65c070df85df8fbf0cc0789;
mem[841] = 144'h029dfd9df30bfe2af93dfe5a0529f002f30e;
mem[842] = 144'hffb4ff050815f541fae5f90f014107bbf152;
mem[843] = 144'hfbabfcf7020a0ea801a10f630337094efcfe;
mem[844] = 144'h02b30729f764fb640bc70c9c0b7a0806026c;
mem[845] = 144'hfd05fdcafc56fb480ad00d6cf85609b9f1c2;
mem[846] = 144'h0cb5f039f2d2fc67f5d200e5f06af2660bba;
mem[847] = 144'h0625fd44f4b20f35ff5e0ed4fb9af6a9065f;
mem[848] = 144'hf0720987fa1a003bf48b0bc00169f023f52d;
mem[849] = 144'hfa2bf83701680f6b0de8fc5e034004080c28;
mem[850] = 144'hfdd5025ef53bf58501f505eb08390dab04d7;
mem[851] = 144'hf42c0c8b00df08eb0ece05b8f4bffa2801dc;
mem[852] = 144'h0959f361fdd7042c0b3a0877fe69f4a107bd;
mem[853] = 144'hf6a7fc9c0c170acf09eff0a9041bf329f803;
mem[854] = 144'h0bb70d27f83afefd03a8065b0ef5f2c0f38b;
mem[855] = 144'h060108d901f1055cf485f414f9e0f558fc02;
mem[856] = 144'h033e0c2cf9f90bb601810d0a015109fefea4;
mem[857] = 144'hf03bf190fbf80154057b01c8fe3006e80d38;
mem[858] = 144'h003e0afffcfafb400909015201c40d76fc62;
mem[859] = 144'h0a7c0a7e0cb50f7c0b990d99f4def94702c7;
mem[860] = 144'hfb150dd80757fa7bf87005dcfda809ecffdb;
mem[861] = 144'h008ffe8800e3086cfe1c0db6fae409fff77c;
mem[862] = 144'h0117fbf2fd310207006300710631027e09e5;
mem[863] = 144'hfd0903e00d4fef6a0856f1530055fd3ff6b3;
mem[864] = 144'hfeed0bc901d6f6f8fc52fb00000b01bcfaf3;
mem[865] = 144'hff51f776026efeeff3dbf5b6fe5609b20037;
mem[866] = 144'hf9dc099af47d0dabfe2df32bf6d3f19b0e69;
mem[867] = 144'hfb82f6f1042308fdf5c9043d0e4bf3760001;
mem[868] = 144'hf0ac0504f6a7ee77eda1f53f0b2cf77e03d2;
mem[869] = 144'h0aac013702840b8bf0490e420405f1e7f058;
mem[870] = 144'hf3ab0151f01104a00d7af104019c0ae1fd87;
mem[871] = 144'hf671f4340404f3d20462f740f360fa12060e;
mem[872] = 144'hef10014ef03fe4c5f547095cfcf5ffaa06a7;
mem[873] = 144'hedd9076d0dcff60d0af5ed84f0a30127ef85;
mem[874] = 144'h016fef8f025dfc6702a006c9fe93f343f2db;
mem[875] = 144'hf8740010f22df862ff0ff8520aca08a0fe2b;
mem[876] = 144'hfff2fab1fc6ffd400bbd08e7fca70408f4ea;
mem[877] = 144'h05cc0ef30be6fd7cf203f89e05a100a20864;
mem[878] = 144'h09ee0a86f56cf035f58d0cbf0cacfc9ef6d1;
mem[879] = 144'hffb40bc1f92f0e8bf89eefac04f2fdb20269;
mem[880] = 144'h0c560f1f0bd9ff5e0910f0c7f7d204920c75;
mem[881] = 144'hf8e2068bf247059f0600f6840d2af5ca0125;
mem[882] = 144'hf175fb00f303ff7ff51ff186f917f179fdb9;
mem[883] = 144'hf2d8087efb900555f7ba0b2106740b550172;
mem[884] = 144'hf0130ac20479f1a0f4cdf1b3f36d0c0defd3;
mem[885] = 144'h035700610c6900b20a3c023bef8ef5b7ffc5;
mem[886] = 144'hfc6202c203def7f70411fb78f9d4f30d05a8;
mem[887] = 144'hf9af0a06f7d7efcaf50cfccffcf2ef65fac5;
mem[888] = 144'hfeabf9acf6be04af07f30140079dfd6dfaf9;
mem[889] = 144'h0b56feff0aa3fd25febaf71ffdc4006e05c6;
mem[890] = 144'hf971070ff712064af27f0d6bfbbe0cb4f510;
mem[891] = 144'h0eba0d90f4c1025c06cbf7520221f933f0db;
mem[892] = 144'hf84cef32008bf06b0e9c0debfd2901c0fe9f;
mem[893] = 144'h03820eebf7c502d00e63f6af0e75fc8e0ee5;
mem[894] = 144'h0b61060b0f8dfbf7f20bf4ce06befcd0f7bf;
mem[895] = 144'h0601f9e70000f4430adbf2730872fa9cfb07;
mem[896] = 144'hf3a1f3cefbe40b31fcb50cf6f16c0285003d;
mem[897] = 144'hf50b050b0268ff46f28102fbf0140805fe20;
mem[898] = 144'hf9eafb1d034f0974067b0bd1f0b20f3009b0;
mem[899] = 144'hf5d1ff80f9aef87cfeeefae20863fae50283;
mem[900] = 144'h072b0bfcf696ef9e0272f195f357f0e000a0;
mem[901] = 144'hf0d8f31afff3f54afbcc030705f9f87c00da;
mem[902] = 144'h08acfb1305560581f4dd024909be045afd32;
mem[903] = 144'hffc6fec90c9905cc04b606e0fee6fb4df949;
mem[904] = 144'hfb1b01a7f2b209e708780e28035cfe2bfee2;
mem[905] = 144'hf7d5081d0056020bffc6047e098c0923f742;
mem[906] = 144'hf784f51909210a83072f0349f282f8af09fd;
mem[907] = 144'h0c9b04ea080ff2ed016f0de407d30df4f4c1;
mem[908] = 144'h0acaf1d408affd4af011fc91f74101fefa07;
mem[909] = 144'hff44f7c908eff028f622012a0759f242f3f9;
mem[910] = 144'h0093f00ff84d09790f3f0b3ffb4c06c2ffc4;
mem[911] = 144'h003afa6a0e6002a30dfb08e1f1540422fd66;
mem[912] = 144'hfe29008608440719080fff0b0ae60cdb0d07;
mem[913] = 144'hfca7f3d00cb407daf34202fb004ff706f5bb;
mem[914] = 144'hfda4f138fd1ef5dd015d04dcf9420071097c;
mem[915] = 144'h039b096d09cd0086f947fa6df5a3fc66f3dd;
mem[916] = 144'h0540eff4fcabf39afefb011dfc6af840f3a4;
mem[917] = 144'h0616ff46f80905430192f8adfeb5082c096d;
mem[918] = 144'h0aacfa29fcc8f877f761fab8ff3ffab2fb1c;
mem[919] = 144'hefb2ef0407f706f30028ff4f0cb3f7e1f5d9;
mem[920] = 144'hf7be0188edcdff8efd0ef7790745efb6faa8;
mem[921] = 144'hfc8fefa403e5fe06f489fddcfd1df7a2f65d;
mem[922] = 144'h06e5f53afe66f420f00ffd5f02e0f7aaefd5;
mem[923] = 144'h0d58f5700479f33cf7cf0d3603daf3d2ff2e;
mem[924] = 144'h000ff34200ccf790f82e08f9f012fa070515;
mem[925] = 144'h0207034a0d8a0718fa27f929f6fc0a960534;
mem[926] = 144'h0641f8b6fddef83bf7baf662f54af10ff736;
mem[927] = 144'h022b0f08fa45f3c802f4f4a40cacf6050a20;
mem[928] = 144'h05160a31f52ff5daf9350d1ff1740427f2b8;
mem[929] = 144'hf918f403fea2f685f402f56df491fd38f7d8;
mem[930] = 144'h03abfc71f803f70ef8220388fb4809200f89;
mem[931] = 144'h0da5f9dbf3280133064cf8fdf7920cd0f05b;
mem[932] = 144'h0299092bf0d3f903fd0bfaa5062609c30ec6;
mem[933] = 144'hfce3ff16f669fa1cef6e0c30f1e7f965026a;
mem[934] = 144'h0020f0550c0f0b500dd4f7e803d8f9d6f5f7;
mem[935] = 144'h0869f3600c5bf0f3f318fd1c0485f8e50a6e;
mem[936] = 144'h0c3df894f44e00ea0e06fb590892f115f6c5;
mem[937] = 144'hfac2033dfc16fe730e4dff6b0d2407f40c60;
mem[938] = 144'h0870fa3ff2d10d5b0d68f1ad0229f7aff0da;
mem[939] = 144'h07c3fd590ee607f109040fe80a280b4307dc;
mem[940] = 144'hf2d5ef3c0e3af76bef6d08a80caaf6440179;
mem[941] = 144'hfceb0942fa98f80e073909a40be7f548fbb3;
mem[942] = 144'hfe2dfb7509d20c1df7e4fb4d0bc3f59cf824;
mem[943] = 144'hff2e02f50f65efa404dbfb0602b40a11f43d;
mem[944] = 144'hf96e0461008ef4ee0476fa7bfa1f00bb0fb8;
mem[945] = 144'hf7c7f279fca1f7c900590dc90026093ff911;
mem[946] = 144'hf7c60baff66b0b31fc94fd8004c3f9daf6c7;
mem[947] = 144'h079f0046f6cbff5c023df0490ceefca9fcfe;
mem[948] = 144'h0d65f5860297f025f2ad09750c540bd8ffad;
mem[949] = 144'hf754fd5cf99bf59d090dfdf7fe5d01fb0017;
mem[950] = 144'h0fe7fd39ff55fde9ffb401f5f6b30b2bf616;
mem[951] = 144'hf0d5f0ebfc8f0785013800060753f075fbee;
mem[952] = 144'h0958fb52f725fe8701230891f022f4f4f879;
mem[953] = 144'hf708fac0f47e0a2801420dc5f77e0628f919;
mem[954] = 144'h0948f6a20afc05a1f7480e8df644f5ba0890;
mem[955] = 144'h0a67f3870773f561ff6f0547035606b8f07e;
mem[956] = 144'hf42ef639f657fdc8f6fcf009078cfb02036a;
mem[957] = 144'hf6a3f7c0f69ff887f0c70799f5e8ff29f69d;
mem[958] = 144'h0e69fd85fd2bf8a70a8ff15cf4eb0cf5f792;
mem[959] = 144'hfb830c53f0b9f6a6f88afa870698f43cfac3;
mem[960] = 144'h0e670e5a0389fbd10c0905fb08fef7b7f262;
mem[961] = 144'h048b0749f2f6f2bbff18f1880225fc9b00ae;
mem[962] = 144'h0b06f0aff5fbffc9f7d1001e035ef37bfa82;
mem[963] = 144'hf02a09c2fe15f45e06b0f87c073dfe4ff819;
mem[964] = 144'hf527f038ef8b0683f21ef06df123081fffbe;
mem[965] = 144'h04d502e2fb04fcbcfeedf76bfb68036900e8;
mem[966] = 144'h052f0d8fff560cbfff8709bbf0f9016ff672;
mem[967] = 144'h01b0092ffae5080bfbfff02c0568f65ff3e0;
mem[968] = 144'hf3c0f7d3f258f0b10ca30dd006a5f9fc08d6;
mem[969] = 144'h0c490bfc0814fae60f3c03490e0ceff4f853;
mem[970] = 144'h0721efae016400f903d7fb7f0362094bf95e;
mem[971] = 144'hfe9af237f1b2f5f2005701c706b008480939;
mem[972] = 144'h084c0d1c0ce606d10aa4febcffa1fad6f759;
mem[973] = 144'hf341fe43fbe103ef05920eb00bc504a60397;
mem[974] = 144'hfb2a066afe4df0690b1cf4cd0a1e0298f271;
mem[975] = 144'h0eb9fafa0a9d0077f119091df3e1f1b10821;
mem[976] = 144'h06350e2f069d0ad6f647f0890f18f199f9ee;
mem[977] = 144'h0e9b01bf04c70684fe0ff665048bf16d01e5;
mem[978] = 144'h0c3cf5760bde0f24029ff53f0830ff7f07f7;
mem[979] = 144'hfe8207e8fbdffa0cf24b0aae0bf10c4a0598;
mem[980] = 144'h0f0cf50b036cfcda0b7b030ff94df098068d;
mem[981] = 144'h026df24e0f4a08f5fa41f1170db3fa18fda4;
mem[982] = 144'hf2f4fa620c970ccd00e00dacf2d8ff2ff325;
mem[983] = 144'h008af7cb03a30850fa04fda305e7f56e08ed;
mem[984] = 144'hf539fe4806ce0354f8c604b303970d56f9cf;
mem[985] = 144'h05ab0a1c061c0843fbfc0bc8ff510cfeff2a;
mem[986] = 144'hf17105250b810d00040af3bffa9700f20327;
mem[987] = 144'h04b2fe9b02abf54c0dba0b2e0ea9f2b2f847;
mem[988] = 144'h0e36f602f2d1fc59015fefd7f03df2b703a9;
mem[989] = 144'hfddbfb26f89e01ae0ad6017ff65ef210fa35;
mem[990] = 144'h0f70fc1efc25fc47f0ebf75f04befdd5f39e;
mem[991] = 144'h0939fb870ba5fd580bb70a7e034bf328062e;
mem[992] = 144'hf6880e47f8c30547ff4f006402ab06ef07c3;
mem[993] = 144'hf5eb0a5c0f350afd096b0035f69bf663fccd;
mem[994] = 144'h0d8f09800352f559f1b0f2fb0c21fc6b07e9;
mem[995] = 144'h019f0b0e07e70aacf9a6f481f7d204180e26;
mem[996] = 144'hf666fecdef61f698f8b2f9c60dcdee8400c6;
mem[997] = 144'h078ef527f1f9f664ff8ff334f6db0d69f508;
mem[998] = 144'h05edf8faf97c0c6f0c9f0aa102a403030331;
mem[999] = 144'h09d506a10926063dfe810386035bf31efcdb;
mem[1000] = 144'heed4f48501f7f0bf082cf1bb0964fdf5f7eb;
mem[1001] = 144'hf26cf380f552f43aee660a840af9fbdf01e2;
mem[1002] = 144'hf856fd1bf2f1fc5b03c20555fa0d038ff20c;
mem[1003] = 144'hfb2cf1c20b550205fc020747076dfbcefdae;
mem[1004] = 144'h047aff12f274f5adf41606e8078bfbb2feb1;
mem[1005] = 144'h047b0a9904d0f3d6f5d20f6bff8ef7c803b6;
mem[1006] = 144'h022c0c66084b0110fe5009d504e8f3bf0d24;
mem[1007] = 144'hf4a8fd77feb60a81f75a052908a9ffd1f0ac;
mem[1008] = 144'h01bcf20df8670420f381fa9a08d5f52c02f0;
mem[1009] = 144'h0d1af36505b2093c00ea0849fad7f1590cf5;
mem[1010] = 144'h01f4f06303aa0e43033e05ee0c9b0d0d0e67;
mem[1011] = 144'hfb8301a6fef1f7a90d47017e0aec04acf6e5;
mem[1012] = 144'hf12007c9fed1f119ee37efa608320c9f09ae;
mem[1013] = 144'hf995fa68096603b50886ff0d088905ed08eb;
mem[1014] = 144'h0370f462f8e50080ff720cfc043cf8160ebd;
mem[1015] = 144'hf206ef4505a7ff21075ffe68067201c8f4e8;
mem[1016] = 144'h0ccf0895fe790d23fe65079cf3bdefa40c32;
mem[1017] = 144'h04d3f578fc380818fc31fddd060eef45f057;
mem[1018] = 144'h0481fcde0cde0363f527f64efc65f43b0b13;
mem[1019] = 144'hf13403e5fd120180f4f9f7bffc64ff64f5fc;
mem[1020] = 144'hfc62fe4402ebfab5f552f858f8e7f30801b8;
mem[1021] = 144'h034b0c6df3fc0c33f0b6fd7bf47cf53ff0b9;
mem[1022] = 144'hfb7c0439f824f552f2f7ff50faf906c7f4fd;
mem[1023] = 144'hf3f1fe33078706ff04f300ec08fff8a9f3ac;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule