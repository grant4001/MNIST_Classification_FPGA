`timescale 1ns/1ns

module wt_mem7 #(parameter ADDR_WIDTH = 7, DATA_WIDTH = 144, DEPTH = 76) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h0673fbb4ef3f02d9ea60ffe4fc95e440e873;
mem[1] = 144'h05ef11950e63131ffd730218fa830390f994;
mem[2] = 144'hf8ccf169f226fd37f60305ecfdf6fa39ee91;
mem[3] = 144'hefb2faa9fe16eb5df98ffe0900aa06540568;
mem[4] = 144'hfb18f5cee636fb51f68409afef9be82ceefa;
mem[5] = 144'he632f1a310cce616faab07d3ebc0fbaa123e;
mem[6] = 144'hf908f23cf95806b5fd6b061205f7fcc8f3b6;
mem[7] = 144'h032d03c8007ef61f07ebf7f3f0edf3ac038f;
mem[8] = 144'hf04eecb7ee31fd280017fa69fffcf5a9f139;
mem[9] = 144'hfbd5f43302ef0197f84f054b0a9ffa15eeed;
mem[10] = 144'he5aef3aae1c90112fb3bf3c4f567e8dbf8ca;
mem[11] = 144'hf19fe51af39afd51e6f4faaaeda6fbe00a44;
mem[12] = 144'h026bed8af4e4f655e9c4013cf759f5350c1c;
mem[13] = 144'h03b10a62ffa9fd1df2d7f89bf5a3013cf16b;
mem[14] = 144'hfe3cf499f5fd08fe012e01bc03e5f4a2fbd1;
mem[15] = 144'h04aaf1c605b1fa8cf86afe62071206e3fafd;
mem[16] = 144'hdef1ff68eccee69fedd7eb0a0074f10fe9e6;
mem[17] = 144'hf3beff77f0e5fc0905e3fc5a1595ffe90437;
mem[18] = 144'hed3d02dbff7bf30bf9fde24ff5ffefdcdf11;
mem[19] = 144'hf57ceb3ae46c00e8f39c0390ffbc0a7ef74e;
mem[20] = 144'hf2e1eeeff738eab5e467ed2be4e9efa9fb9d;
mem[21] = 144'hfe32e5a5eb21f93aeedff797f6beed51095f;
mem[22] = 144'hf791fa4c07d3e7a9ed1701c4f2fdff4bf700;
mem[23] = 144'hf509ea5af661fff8e804f60ef4d5013903a1;
mem[24] = 144'hebdef9b7014c04a0f3caf196f0c3f789f518;
mem[25] = 144'heddcf845f28efe9a04fbffe3fae8f6130185;
mem[26] = 144'hf8acf13df682f85cf23e053100e3f0acf4f6;
mem[27] = 144'h08edf095fbe4edbc07160c18fffff21df7ad;
mem[28] = 144'hf291fce5f880025e098dfe47f6e1f42bf8a8;
mem[29] = 144'h03010247f005f6050198fe79000afb7ffa19;
mem[30] = 144'hf022fd6beec6ed1cf098fe9afea7eac3fb8e;
mem[31] = 144'hed72e9e6feb200a1ead2faece4d0e665f9c1;
mem[32] = 144'hecf5f9f709b7e99e060ef144f4d9ecb90559;
mem[33] = 144'h0954f015f595edbf03b9ffd8f753fbedf7f4;
mem[34] = 144'hfee8ed1df4a8e1c9ea48e884e42ee073ed85;
mem[35] = 144'heb24fac8f0e3f1f8fb3ce9dd0250042c0cf4;
mem[36] = 144'hefadf052fcc8ee37fa5afe70fa6904b80679;
mem[37] = 144'hf5cfec81f552f8a30732083dec7afd52e8e2;
mem[38] = 144'hf6b609c0f32cf8c6f387fd6ffbc3eb5f01ad;
mem[39] = 144'hee5df881fb2dee2df70ee34eea17eaf5e96b;
mem[40] = 144'hedb5f7a6098ffd1705240435ef85f494f9f5;
mem[41] = 144'h08a0fc3ef5e4fa90edfbf4acfd320937fff3;
mem[42] = 144'hf15bf569ece3f2a6eb70fbe2f222062adede;
mem[43] = 144'h01f7ec51fd18e94efb84ecaff0d1089a11f4;
mem[44] = 144'hfc93fadcff98eee605d10855ec7deeacee0b;
mem[45] = 144'h078f064a1b020c3b1f4d276611d713440ff7;
mem[46] = 144'h01d4085df6ccedd1f658ef6ff95800c6f7e6;
mem[47] = 144'h05f6ed3ef6e60991fe15fbb1f8cc03b4f289;
mem[48] = 144'hf6b708be033bf50c052a05c0fdf302a40342;
mem[49] = 144'hf959f793f17dff8205d6013101200536fd43;
mem[50] = 144'heedf0922f710fdb104f202950810f94f0804;
mem[51] = 144'hff63fcb9f632ee27f5feee34f763febb073c;
mem[52] = 144'h029ff8bee727f046f514e9a8f83ae71bfd0f;
mem[53] = 144'hf39af49ce550f39eeefef823073407830305;
mem[54] = 144'h0957efb3069efbd203eaf4ba05fa0936f3f1;
mem[55] = 144'h0775f3b204faf4ac07e0ed280661f1abfffa;
mem[56] = 144'hf3a9f4b908480385ef13f152ef6e09b2fa92;
mem[57] = 144'h020d01bdf755f8f3f8bb0a0e054af661fba6;
mem[58] = 144'hfa2efdf204840867f30309a6fea40b410403;
mem[59] = 144'hf27cfb1bf7f9fe460b53f0a1fc6ffc77f607;
mem[60] = 144'he560e3b0e00afd8cdf32f763e319e96cf666;
mem[61] = 144'h0c8bff2aee1c001416f101acfab1f42c0b6f;
mem[62] = 144'hf05ced130172f160f7a6ecfc04e1f47d05d6;
mem[63] = 144'h055debd90230f3c402f5fd51edd50326060d;
mem[64] = 144'hef4bfdf2fb57f75400f6fe78ea9ce538e19b;
mem[65] = 144'h021bf831f573fe6a0f380853fcc6ee8400c1;
mem[66] = {16'h029f, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[67] = {16'hfeb8, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[68] = {16'hfebb, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[69] = {16'h0509, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[70] = {16'hee59, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[71] = {16'hf137, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[72] = {16'hf5af, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[73] = {16'h02eb, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[74] = {16'h0832, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[75] = {16'hfc29, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule