`timescale 1ns/1ns

module wt_mem3 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'hf9b90d78e2f40a79e20ae61deaf5f1b813fc;
mem[1] = 144'hf593f3eb0623ea6101d4f0c612fbeaae0949;
mem[2] = 144'hf69ae2c10ed4148eead00975e0fc098bfcdc;
mem[3] = 144'he1dfff45fd5e1b7205061da30ebeef3002ff;
mem[4] = 144'hfd0be558f907fbade887153614d2eb19136b;
mem[5] = 144'hf6021a01f0b00561184d060ae6e61457e171;
mem[6] = 144'he24afe4e06dfeb41e9c6ec460e31f5d50f42;
mem[7] = 144'he601171d0af901a0ff080f7101f1f92e0148;
mem[8] = 144'h0c9618421763054c1f4a0733142fe0081f5b;
mem[9] = 144'h07bd1b99e40f04b70ea21711e3550f381bcd;
mem[10] = 144'hec96fd30f541e5fae682f308f3ac1fb5e3f9;
mem[11] = 144'h0645ed30ed2a1285e58cf8d9f78811670350;
mem[12] = 144'hebce1a7cf40fed920d3beaa3e4f303b307d7;
mem[13] = 144'h019af987f058f4dafa91e15002f9eb911b1d;
mem[14] = 144'h140a04d5efe9f88801ecfce80781f19bee93;
mem[15] = 144'hf834ee5afe8f0d14f13807eb0eb00b13ef22;
mem[16] = 144'h0a690d830a45f20407f9e30deebf05cef654;
mem[17] = 144'h02cb15b203e31f07fbbbf1390dcefe1f0ff0;
mem[18] = 144'h10ce0b16fa12187b0a84f19ef23de7dc0dde;
mem[19] = 144'h1b9719770738ec3605f91471f08d003f020a;
mem[20] = 144'h00540081e54ff15f057a0a57e67310d30116;
mem[21] = 144'h0b860359ee980d2eedf5f7bc094a116e1905;
mem[22] = 144'h0af9e3a50bf21594fcd20e0b1e2d0547099a;
mem[23] = 144'h127f1024f146f457e7080194fcf1e7061e40;
mem[24] = 144'hec66e28203c3fbac1c90ebc30ff210dfffdd;
mem[25] = 144'hf3e9e5f31a8fe48ffdaa0922eba5e099e017;
mem[26] = 144'h199bf629146bec62facb07ff1048e9f70f44;
mem[27] = 144'h1b7d029ef4dafa36ed4ce624e006ee090fd8;
mem[28] = 144'h075814f1fe731f6f0b41f98aed09efef065e;
mem[29] = 144'he6f0044c0a66e2501d91017e078f0fc0f0a2;
mem[30] = 144'h09a3182aeb840e81e0eb1b48e60cf2d6e45d;
mem[31] = 144'h0278e255f75df210f4e1f3c91e761e46e7bd;
mem[32] = 144'h1b5f05dd1319e464ed03001cf32a08b209a7;
mem[33] = 144'h148b195706d008d300fc10abe10802d916be;
mem[34] = 144'heccaea6410f206dfe05dfaf302c11160e3a3;
mem[35] = 144'heeb018db0d8de57aeeec17dce45017241c08;
mem[36] = 144'h1439e1c5018be64b198ce7b117041999eb61;
mem[37] = 144'h1e01095e1a5d14c5f84be0f31d6afe80ea07;
mem[38] = 144'hee81e45efa3a023ae570e7e5f286e45ffc5a;
mem[39] = 144'h1b0df59ff7f0041d0e201b0dfb9de0e002fa;
mem[40] = 144'h0201e911fea0133efc0705980f49f66de955;
mem[41] = 144'h1c8c00a4e4f6e5dc075b16711a24f43be940;
mem[42] = 144'h1bfff0a3f6d500db1093102fef6b1f93e70b;
mem[43] = 144'h1e7c1defe01e05f819580d8ef37bec291789;
mem[44] = 144'he238fe51f8bdfcdf1ce1fb9de0e2efef152d;
mem[45] = 144'he47af25500c61ccd0bfa0e2aea20e9091b72;
mem[46] = 144'h045ef73cfdf8f85dfa130036089bf7971a44;
mem[47] = 144'h02a80bd3f4def206ed52185efec606ebe889;
mem[48] = 144'he6a3ef71fa72f82807deedf0f0d2017716f2;
mem[49] = 144'he393fafd1004e8d8fa531ec8173c1d62eef1;
mem[50] = 144'he292088b1074eef01f1d18baf71ded42fe3a;
mem[51] = 144'hef28162917201612f7b2fdb11442f8870484;
mem[52] = 144'hec0eef971a81e17617991e55fcc301d50578;
mem[53] = 144'hea96edae0012eb9ff3141a340c40112ce3b4;
mem[54] = 144'h02bc161ce7851722184000941a2f0fc2eace;
mem[55] = 144'h02931bba093be6821e2fe459e284f71aed4f;
mem[56] = 144'h1b920a5af6cd1e940694fe70e5fdfe530af3;
mem[57] = 144'h094fe638ebfb00defdad0720141f05c0e353;
mem[58] = 144'hf80ce88a179517420b0c1013f2afecf7fad7;
mem[59] = 144'hef35fdd810fa14531ce604c5f9f91dc21a9e;
mem[60] = 144'h085415c9eb741ee9fe01089b057402e51da1;
mem[61] = 144'hf256162efb8ce4f4f953faa319a3ead40ea4;
mem[62] = 144'h0a35f9080dd8e0d5e2251af70df5f9fc1efa;
mem[63] = 144'h0b7eff6ee4430457f980fa4e09b7fe8f1e06;
mem[64] = 144'h103a0234066f1581fbda1c00f03dea1be6e7;
mem[65] = 144'h1a2e0800edb519410454e040f9811940185c;
mem[66] = 144'h11cbe9a01abdfe791345e294faa50ba30c92;
mem[67] = 144'h18ddf84f00bc1252f66b1d77ef58fd221cc9;
mem[68] = 144'hf2e505abead4119700f9f266efe90c14078d;
mem[69] = 144'h119ef3761b3a09c202bf058d1050f9431f98;
mem[70] = 144'hf6ce13ff1c67f66c1802e686fd5ef2340439;
mem[71] = 144'he450f880e52e18aff77ee56909dff3def35c;
mem[72] = 144'he77a1183eddce9f4e861062cef2e150fef3c;
mem[73] = 144'h168615caf33eecc4126cf1c216e9ebb6f6f9;
mem[74] = 144'h05b317c1eef00537055f09860e88fc61e31e;
mem[75] = 144'hfc08fe0e18d6e75c1e7afa5afbdeed50e3a4;
mem[76] = 144'hf009e2cb00601a21f753e013f124eabd115f;
mem[77] = 144'h082bf2a1e24810d8180ae2680432e54af633;
mem[78] = 144'hfd85efa3160f172a1dad060c09d8f5241f57;
mem[79] = 144'hf1cb0797078be2580768e52de865e62ae8a4;
mem[80] = 144'hefa30cbe06eb021c0e52e9f1f78be0eee247;
mem[81] = 144'hec78180ff5241d0d0d3a06ccf0b91f29f39e;
mem[82] = 144'hfb4ff55bfb801fadf32d004d0f5909a6e619;
mem[83] = 144'h0c5c10f3f515067d182df14609d4070fe0aa;
mem[84] = 144'h020cea68f18d009404f31783f075efbfe494;
mem[85] = 144'hfd1b1c8f0b04034df49ef44516441930f426;
mem[86] = 144'h1f49ece40bccfd7ee378f7ac17661448f45e;
mem[87] = 144'h00991f4de499e1cae251fe96ec80fb4c0179;
mem[88] = 144'hf10000121c75f38ee7d216c2e8f6fc0e188a;
mem[89] = 144'hf8e6f8f3f8610886070c1e0ef92fee5afd6a;
mem[90] = 144'h018d10f5015dfbdc0d180772e20ef52c0feb;
mem[91] = 144'he95c1cd6e72f1e4f1ad81cd4f46e0512e4b7;
mem[92] = 144'h0ff51e720812107df2ba00fde837156b09ee;
mem[93] = 144'h01e4ff31e0c2eed5eca911a3eb2afa14ebc7;
mem[94] = 144'he338e6691dcdf577ef2ee90e1dc40c2aecf3;
mem[95] = 144'h032a000fe3ad1635fe26e159e72e0330f0b2;
mem[96] = 144'h0a731d65fe4d1291ea2eea7f1829f0b91bcd;
mem[97] = 144'hfdd9f93bfa91110fe48afceffe4cf91607e6;
mem[98] = 144'hf1eb036fe51aff6611a4193f1926ef31efbc;
mem[99] = 144'h1c291ac8e0161c9ce0651cc3f77502d1eabe;
mem[100] = 144'h007ceb44e050e1a6e051170eed6cf108ec0f;
mem[101] = 144'heea0114ffb1c011defb30d68ea5dfe12e295;
mem[102] = 144'hfe420df70b5ffa62e4b000b511d405db1f8f;
mem[103] = 144'h034407dee1800855f2cd119a11c4f87707fe;
mem[104] = 144'h0fe3f536023d0f2ef5e3e6da1391e383e20b;
mem[105] = 144'h0ba907e3066de71e04a0f1280c541d2cf08c;
mem[106] = 144'h0fc1ff9ef8680d1700a7edfa0275e990019a;
mem[107] = 144'h05690042171e144de0f21b2e07ba157e17b3;
mem[108] = 144'hf60af9c0ff8ce4d71587ef760433027b0f47;
mem[109] = 144'hfae81838ec8e169604e81b61fd01f04d19a9;
mem[110] = 144'he53cfb531c08e574fc0417221ccb0022fefe;
mem[111] = 144'h096703530319fe3409010b0e1ebdf6c21a8b;
mem[112] = 144'hf3410ce80c8e1cc81ba3e9f0e5451da21007;
mem[113] = 144'h0e26f121e04315a1017cf471eed317d8eee1;
mem[114] = 144'hf5580338049e00390361f8b0e1a8fe8e1bd1;
mem[115] = 144'hfaaf0c59052a08660c9319befece012e1056;
mem[116] = 144'hfff20fd8f9721e6ff68b033e0529e874f57a;
mem[117] = 144'h1bd014adf472f9e9e169e48dfb3e075cf622;
mem[118] = 144'h1c050c26f8451c9cec59f4b6f5d9f916e1ba;
mem[119] = 144'hf3f4fa0304c9eed7163de97ce43007ece041;
mem[120] = 144'h06d5155315d40677f8e503851381ee1c0ead;
mem[121] = 144'hfdec1435ee7f1e1fe060f9d21ebee868f5ff;
mem[122] = 144'he944066cf1fc09ab04e21f29021817f5ee8f;
mem[123] = 144'h1f920cc3ecf406f408121d6d0cece299176b;
mem[124] = 144'h0e2ffa26f5371ab7eb8ce01c1e7a0c09fe2d;
mem[125] = 144'h0ad8ef32f73cfe76f9a2095affcf100f04ef;
mem[126] = 144'h105e04470727120ef3260c6f10511aa8e320;
mem[127] = 144'he2f000f8047bee5ceae91ec1e632f2c10510;
mem[128] = 144'hf848e9af0b61ec91014419431509e9ec0571;
mem[129] = 144'h01fd0c95e9781601e467e563e974e998e4af;
mem[130] = 144'hf77cea45153c11340380f2b1e8ce1beffeb5;
mem[131] = 144'h14411e33eb03183ff5a3ec77f9bbf255155e;
mem[132] = 144'h1a561c80e1b3ef8302ddfd441573f608f3e8;
mem[133] = 144'h080be7741f7b029deb0fe5f7134be87e1523;
mem[134] = 144'he780ead1178f1cb5032919a20fdae76cf180;
mem[135] = 144'hf7b1eef1f4cf0dc0feb0f3abe206124d11af;
mem[136] = 144'hf6000ee01de905e7f15ff3960b141890f284;
mem[137] = 144'he9bb1d5503761c7f06bdf1451adbf6801999;
mem[138] = 144'h130ee40e021ee7ff1dcf0c42e4ce04c5132c;
mem[139] = 144'he5c61285fc07f2271d7bf459e8c6ed290926;
mem[140] = 144'h113f0f4ee02a0dce1424f8a4e3fa0f7701ac;
mem[141] = 144'hf2df0e17e9790963fad00885fa9d1f2eee9a;
mem[142] = 144'h09e0fc6d1adc02921de5f9c0e406ee55f914;
mem[143] = 144'h1bd206e4e2f8e1dafcff16d206a0f842e2d9;
mem[144] = 144'hec56fc740ab9f83ef393e90afa3f1813090c;
mem[145] = 144'hf90df71dfd4b1f8e05111b54ee86fbf71bc5;
mem[146] = 144'h12dee77ef63bf8d60ec3eefafb24ef6e187b;
mem[147] = 144'h1383e813ec79e7daf3850ef9f55d184206c6;
mem[148] = 144'h0ebe0a1c16b319aae5e4166716921048fae5;
mem[149] = 144'h0eefed031048f1841cdcebd3ed361575149a;
mem[150] = 144'hf472162903bffd7802f70cee07fd1fc50026;
mem[151] = 144'h0ff31dcd0198e4db00d11f081fe1060eed98;
mem[152] = 144'hf66ce23e1f441a5be24b1bf7fac4042506c6;
mem[153] = 144'hef63ffb9f4bc0935efe311f200fd1aec16e6;
mem[154] = 144'hea7bedcf08cff9fde97008921f0b1facf4bd;
mem[155] = 144'h05f4e8d31f570ece197500a81eea02060951;
mem[156] = 144'h1f9cefc715bd0b4813f0e54a104902f4f671;
mem[157] = 144'he391f3dfea72efb3ec1704ad155bf13ce09f;
mem[158] = 144'h0587fb060fb4047df573140908a2e79df4d6;
mem[159] = 144'heaabe38d072ce692f782efec15000400ef9c;
mem[160] = 144'h1ed905830f30163c18e3ed651b83f7bdebd7;
mem[161] = 144'h0f7610dbe583119610b5fb351c55f318f18f;
mem[162] = 144'he27af98211eafd021183ecdc10efed6211e0;
mem[163] = 144'hf710095fe99e1411097aeb31f1201bf00125;
mem[164] = 144'h199502ceed1dfcb2f16ef642093618e9e59e;
mem[165] = 144'h158705ecf4d3e9eff5a8ec520a09fc97f4f9;
mem[166] = 144'hf926fe38f335f7b1f0c2e7a10e7ce031f7a8;
mem[167] = 144'h134fe945f9b91e1aedb4f94d0c5709aced0e;
mem[168] = 144'hfe691306f7910049f86ffac6f6fcec4e116c;
mem[169] = 144'hedf715fd0dcffb6df3ba0d76088ef9530517;
mem[170] = 144'hee03eabcece7e0bd11a0fb49e207f11313d8;
mem[171] = 144'h1e61f4450a65e20a11eee3b71f9e02baf67d;
mem[172] = 144'hf45fef90fe3a02730da300abf35f04b91b97;
mem[173] = 144'he8400d4fe3f40d340ca3079a0583fa2d0956;
mem[174] = 144'h1d1f11ccfcb1088bfeb413d5fc5e01220989;
mem[175] = 144'hf728f33e058be5591ac3f56fe3960fe50ef4;
mem[176] = 144'he319f1bfebd2084e11a80244f29cf182ec47;
mem[177] = 144'hf97df53be3e1f906190b0241e961181fe77e;
mem[178] = 144'h0e8215350d55e88119a7f8570190f170e12c;
mem[179] = 144'h1a7cf8b900591e911af4e6bb112313991c58;
mem[180] = 144'h138406401710e40505ceef431f0a0d7803d5;
mem[181] = 144'h0615e084f836187affe7ea2bf2ac1af31aab;
mem[182] = 144'h14de0d8e1636f58ced641fd80afbf00dee2b;
mem[183] = 144'h0631f9990854f9e51b390aaf1cde05c412de;
mem[184] = 144'hf6e51050019412b403eee1c6e756e4fc1cb0;
mem[185] = 144'h053802e9eb2615870d2b109df862182fe220;
mem[186] = 144'he13ce316fd9aebdf0c2215ca0b02eeb11fe7;
mem[187] = 144'h19951b97ec180fd3fb6407d110ca1f62e445;
mem[188] = 144'hfe5507bc1cd21f5a1c9f01bce39ef9d6fdc5;
mem[189] = 144'h09a4e3d9f6e707a00d1be52bfcecee0e0e53;
mem[190] = 144'hec171bf6e66bef82fd830286031c0492f862;
mem[191] = 144'hf1e814a2e7a50ba7046901daecd50888001b;
mem[192] = 144'hf261e8b8f311f4bf072210a2f4220b680103;
mem[193] = 144'hf254f7e2f275e95d18dfef8c007bf5cff244;
mem[194] = 144'h17daebd705d2108be8d80611104911a71154;
mem[195] = 144'hf27403fde11deecd1928f41aef621e050f70;
mem[196] = 144'hfcabef04e398e65ae04ce3431ea8efc60aba;
mem[197] = 144'hf944f1650461ec08f7b1f16e0be4114e0845;
mem[198] = 144'hea39f2f7122eff420f1d1c64ff060ae1f8ba;
mem[199] = 144'hf2f2020d086c152aea98116618d3ea2ff146;
mem[200] = 144'h0ea70c5809b61380f2afef12e5aeec21f055;
mem[201] = 144'hf4ae068219bce941ff9fef04e5cf0666f173;
mem[202] = 144'h104f02a3e6c0110ee7911d40fa27005b17cb;
mem[203] = 144'hf1790e921eba1c430db8f09bf6971fb7f4a3;
mem[204] = 144'hed3c18a50588e7f710c51935ff19f6540336;
mem[205] = 144'hf63f1d4d1f1c1c2f1908ebc4f03f1284f3fa;
mem[206] = 144'he0b8f770f87104ed0e4ce51cf22c03270bfd;
mem[207] = 144'h0b08f9100dd00319e677fd81065b13a50ef4;
mem[208] = 144'h1ca50cf1f4500e0f110cf8a51e4e195304d2;
mem[209] = 144'h1219e9c9e854f1a70aa5037a0151fc04e14f;
mem[210] = 144'hf24b000df820042d12d2f12deadef5350be4;
mem[211] = 144'hea89ecaafe261a6a1fd2f6521d8201890cde;
mem[212] = 144'hef0a1477ee4ef795e1f8e8a30bb0fce4e761;
mem[213] = 144'h07840a390edafbe40a4beba1f3b0edbce498;
mem[214] = 144'hee9dee5a1e18167ef9f2122e048907aa1378;
mem[215] = 144'h0b5ce675f5edf24bf24a073f1d84e2ad152c;
mem[216] = 144'hff4fffe3e9c609a8e1500fcdebee1db7fa8a;
mem[217] = 144'he19afc57e3d9ea9f1dd9fb45eec001811041;
mem[218] = 144'hfa881cbef6a5e8f810941d35f6c0fc8af504;
mem[219] = 144'h093f17c6033a018fe4bdf3ec0db6f0e01d71;
mem[220] = 144'h1235ef3ef0b7191a099cfba61ed2ec2be06e;
mem[221] = 144'h100dfe670eebeae2ea3df668fb3a02060528;
mem[222] = 144'h0ed4f7c4ea6410ad15f91afcfcea08ecf464;
mem[223] = 144'he103f37beef3020b041907860b93fb2be2b6;
mem[224] = 144'h079ae7b71699e9baf96b072febcbe0c00b96;
mem[225] = 144'hef2f16cbff900ec9fa6a0f0b01adf75e01fa;
mem[226] = 144'h0a0ae816f9340983ec1f07d60b0e06991788;
mem[227] = 144'hfd2df936e2f30b4ae4aaf9891b1be7390fa9;
mem[228] = 144'he44c1277e2e600def81c050012451b99f434;
mem[229] = 144'h0b57ecd9fa3df73cfdcee2421c55e90b0b70;
mem[230] = 144'hea7c19c31e9ce45d00fe07cb133afb021237;
mem[231] = 144'hf99d052b1d3ae0f6e042eb64e671e8c51fd3;
mem[232] = 144'he3b8ec77e59e0657f1cc19471ac8f842e19a;
mem[233] = 144'h06990ba513411a87e34ce9e7e562e5eb11d8;
mem[234] = 144'hf9b0f2a60ac2fc9ef558ff8df073057709ca;
mem[235] = 144'he867e5cefc8d0a8b0646e5d5120bf383142b;
mem[236] = 144'hf876f566e457e19b052802f0068b1213f38a;
mem[237] = 144'hf2dcee680edb0ab0f102e7a0e2e5f3d81ff7;
mem[238] = 144'h09571088f68c01d5ff300e1d00d6f0a9e6f6;
mem[239] = 144'he4cffe4c0fd4edabf4d10b5c0e77f863f9b2;
mem[240] = 144'hf975f1b4174719840ab9e364e8f4fcc5f5c5;
mem[241] = 144'h1f19f744e0e2e6e9f8481b97fa2be09eefe6;
mem[242] = 144'heed71756fb691313e1db137e0798ebc70527;
mem[243] = 144'hef8af5c7fc4e0e67e84cf22cf18d099d17ed;
mem[244] = 144'hf23005b31010f853ea9819e1f65307671ec5;
mem[245] = 144'he11c0be3074618631922e48bef4ae73bf700;
mem[246] = 144'h04590780069c01ae0d7a1cd8fcbe085209f2;
mem[247] = 144'h02fbe6b0f55604defbebe14019a2f217f94e;
mem[248] = 144'h1ef00a8cefd1f31208010ec5119c0ed3fe05;
mem[249] = 144'h02f70b10e0a0fed01b57e1231f391d340bc7;
mem[250] = 144'h13ecfe9ffe19f6f00b4f11b2f2cb15a9f032;
mem[251] = 144'h0e76f4e00bca046d0871e91c14eff40efe75;
mem[252] = 144'hef0d05fee52bfc3ff26f05be147209c4031f;
mem[253] = 144'hed6dffdb131e03effadc1750ed690a56e316;
mem[254] = 144'heab7e52909fee2baeec7eb25ee0a0040185b;
mem[255] = 144'he62ffad7fb0e049813d7ed50f8300240f633;
mem[256] = 144'hec131f69fb911578f0b6fbd4ec67eb35f453;
mem[257] = 144'h0b88f29ef508e59205aa16f3ea17e9a61ed2;
mem[258] = 144'h07ce1111fb13ee1ce827e6a7e070e5990812;
mem[259] = 144'he01ff6d0ea780be41ed2f417ee4aec371db4;
mem[260] = 144'hfba2fbec0cade01cf399115b11f4f08818b2;
mem[261] = 144'h0f4be6d11e331348f09ce16e0cb4ee5ee9d3;
mem[262] = 144'he9aceea9e0e2f50b1f70e70ff186e266f6e0;
mem[263] = 144'h095606230af2e3aff899eca101e1106d1994;
mem[264] = 144'he49eea70e8cd1dcfef3af2581641e7cb0853;
mem[265] = 144'h06be1ac3e495f98cf10903d5fd8a0268162d;
mem[266] = 144'he23cf01debfcf422f974f67cf199f9721b74;
mem[267] = 144'hfbefec8d00f317a4f870e99a0267089b1e52;
mem[268] = 144'hfc49e4b20a72e0d0e2761b88fad0fe3ff0fa;
mem[269] = 144'hf2c9f9c31444054e1ce1fa11ef04e6e0f1e7;
mem[270] = 144'he4a813f8f9f1f0dafe4be0d712eee4f11c00;
mem[271] = 144'h1874f717085b1f330df10110189c183af377;
mem[272] = 144'he804e7261e6f02120647f0a9e7d3f26a1b22;
mem[273] = 144'h049b1c6f0a18e982f3be16fc0aebf872eda2;
mem[274] = 144'he4cf041eee0316e8e88f0eac0f60f3c5e71d;
mem[275] = 144'h0761f7dc048f12fde5c70df8f02216d51ed7;
mem[276] = 144'hfd21032f1acd0dedf1470d11e2f80864e175;
mem[277] = 144'he348fc53166fe0610b5d06d7e8baee35e32d;
mem[278] = 144'h0b1c0509efedf5e5e9ce17900e03fc50f5b4;
mem[279] = 144'h0c36fe63e15106a61f4a02ba13d4fa3001f3;
mem[280] = 144'hf92ef8900da91b08eb8012601f6706e80917;
mem[281] = 144'hfed806c4f69401381c10f93610da13e30956;
mem[282] = 144'h0be5f47ee1e6fca5e88b191aefda1339fc29;
mem[283] = 144'h021dfd601082f2f6ffadf3dfebbfeff8ee31;
mem[284] = 144'he20e0df811a60c0ae903e931165507e507ca;
mem[285] = 144'h026b10040960e5350dc114b5e1ecec7af76b;
mem[286] = 144'hfd4e11e511aef4f8013ee6e3eb04ee541581;
mem[287] = 144'he4d2f078f7c0f29b148d1d8fe944e330101b;
mem[288] = 144'h0d3df5d7110ff200f947000c0072f711f70b;
mem[289] = 144'he2c0f8930054f9060bae102a1e6a163cefde;
mem[290] = 144'h1ddff8efffcb19e7e83609821f79eec7edad;
mem[291] = 144'h0a51e762145f01e50bea1c75efcf1c581acb;
mem[292] = 144'h1eaef6971a2cf616f3a9fb09f6950c841740;
mem[293] = 144'hef92e81ef89f05bb01fbf150fc76ee331418;
mem[294] = 144'h1974e883f3bf0ec9fe531113f950f4eee35e;
mem[295] = 144'h09f8143e17270780f0d2f3d61001e94ce543;
mem[296] = 144'h0f6fe9c6e0d5099e11a7ee7e0fd2ef210034;
mem[297] = 144'h1fc8eed9f9e81ab00932eb6e0fd202b2101d;
mem[298] = 144'hf0400740018f1ef607770898f372f250010e;
mem[299] = 144'he7e8ed3b0e0ae0aff9831709f139ff5bed1b;
mem[300] = 144'h151bf833eca609a9fd5be173e907e0371f53;
mem[301] = 144'hff040574e694f0f4e837f7a6f183e982f6e7;
mem[302] = 144'he0d7ee25e6e206c4e7440cf20bda0bf01bc1;
mem[303] = 144'he15eeed20a7216a8f4fb15e10f28f6831839;
mem[304] = 144'h0e730aa4f66800bb0f141f54e9cd109cf05d;
mem[305] = 144'he9f718ae1551f8bce0d61843145a0230f1ad;
mem[306] = 144'h070aff5ee28df2b01bdbfe61e8341a30e254;
mem[307] = 144'h0a430018e57a104c1b74e59eef56e6a2f225;
mem[308] = 144'h1b521fbb138e0a0205611d4ef6d9f9d6efae;
mem[309] = 144'h0ebe015bf195fa09e2f1fe0a0954fc8518cc;
mem[310] = 144'h0adde43eee881553fe8f0b9af8de13111727;
mem[311] = 144'hed6a04d6f58f121fed14eceb191a0f13fac9;
mem[312] = 144'h0c81e38e07afeb3f15d102efe37d1216f9dc;
mem[313] = 144'hf3f9e96efbf70aa3fe6c125dfe200ccc0bed;
mem[314] = 144'hf3dd0f21f8930d5d12fa05620f9ee904e6b2;
mem[315] = 144'hf429e952096afb52e01b09bc02d1f77ae8e9;
mem[316] = 144'h182b1ae2fb3d02f0eb4dea8f03a3145518ca;
mem[317] = 144'he3e6fb8901b006d71a571726fe2ef0cbf8b9;
mem[318] = 144'h12f301d31ce1e73dedd91a5a15c5f95d1ee5;
mem[319] = 144'h0726e5b700fdebb6f246ee560322f987f9f9;
mem[320] = 144'h1e570a48f5f10a37f5e6f082ea8afe420d6d;
mem[321] = 144'h0195f92df61f1227e916f57518091369121e;
mem[322] = 144'hf88f18c304260e75f17d1bb5f7141bf6fc73;
mem[323] = 144'h0b8a1440eee5003ae914f1e4fb66f2f6e3c0;
mem[324] = 144'h063ff75c1ffbead60277105be84eec62fbc0;
mem[325] = 144'hfba8f0511560e1fb0b66eb3ae56af3cde0c4;
mem[326] = 144'h095beca60e320d4cfb260e1606a616aee4b8;
mem[327] = 144'h1cb2ed4f1ade02e2e610ffec13e80acbe135;
mem[328] = 144'he0620c221e4deb720a09f51ae12df3a50437;
mem[329] = 144'hf131eafdebfbe6671265f3c7fca11f1be144;
mem[330] = 144'hfef91f72035c1fad05ac0ef4ee530f1b0cc9;
mem[331] = 144'h011e1360e5a1eef80f9110a8098be28005ff;
mem[332] = 144'h1c88082409ce0ce0f4d31a111d7f050417f9;
mem[333] = 144'hfe931d21f1bdfa68ebe2f215eaa015170c86;
mem[334] = 144'h088bf423ed48f5e10afdeb0519a1058df393;
mem[335] = 144'h09c4ecc30a5d00371c59e70df6ecf6f3f613;
mem[336] = 144'hfccb18ab0164f097ecdd12d9f4a0fd6307c3;
mem[337] = 144'h19d6f61af081e754f5981768e927eb54fa46;
mem[338] = 144'he1f519ece325f5b91c55e62cec3be20af4e7;
mem[339] = 144'h1671f5fcefbf1a0d189a062714dc1323148b;
mem[340] = 144'h055b1dd6134007c1129af76d1eddf3a7e8aa;
mem[341] = 144'he018ea3bff81fbacf31813e900c4145deffc;
mem[342] = 144'hfa6feea8098bea1fff3106cce1291b150bd1;
mem[343] = 144'hfe9dfb96efc0fe56e8e406fcee4108ab19b2;
mem[344] = 144'h02d6e45f0586f4d2ee3e0b0413c9f2bf04e3;
mem[345] = 144'hed211031e36f1b74e08701b61371e5c5ef2b;
mem[346] = 144'h14f9e1451c5ee88c0425f65d00ace3e406d3;
mem[347] = 144'h019ffdd205a3fca2f7bfe80f0571f997f1dc;
mem[348] = 144'hf977009f1cc2eea6eba91f0c17fd1d761046;
mem[349] = 144'hf6d1e2a50dbd0302f2abf7941e07e78c0ece;
mem[350] = 144'heedf02b81e6b0911170efc2be557fa45164d;
mem[351] = 144'he2efe1e714820858fb990b1df114fa59f30c;
mem[352] = 144'h1bbbf0ba0d2304f5fb5ff9dff6b7f0f1f24d;
mem[353] = 144'he7ebe688f8820560e330efda17700d9900c3;
mem[354] = 144'h16e2ffe617d3f17408d706580db905fef263;
mem[355] = 144'he263ffe8f686e7e9e14415050780fc45eb7d;
mem[356] = 144'he73de195f4abfb2df7db033dfa9c0c59edcc;
mem[357] = 144'hee6efb0dfe1dfa72e6bee130efed058ee36b;
mem[358] = 144'h0aa609431b5e1e841fa3e8bd0c62f2ce04b0;
mem[359] = 144'hfdc8fbe0e50af5431b8813e0e9f002c5f802;
mem[360] = 144'hf9b20492004f088c05300cbf0bed18b7104a;
mem[361] = 144'h1766e4ee1b87ee7de979f3df06691cc5f509;
mem[362] = 144'hfbdc1a0b03c3e10feb9315cb075f0cc9018e;
mem[363] = 144'h03ec1d51f24102240c48110b0be6075d03d2;
mem[364] = 144'hf6f20b8b0dc5e9ce14eeeffaf26d1d270c59;
mem[365] = 144'he835ed98ee9f10fe08281846f454f04df9a1;
mem[366] = 144'hf61b0c7e004eea07e4c4f2d0090eecd40755;
mem[367] = 144'hebbae3530f9ae599f55e0e7317f407060db3;
mem[368] = 144'h00b7117a116bf4e5f2ba0ef71a98eab90f42;
mem[369] = 144'hf4d91406f901eb360a7517d108f40b9a006c;
mem[370] = 144'h06a001df170beae617d8eef3eb62e2ceffc6;
mem[371] = 144'h0b92e78efa2e168bf5ef120fec68ff85e23c;
mem[372] = 144'hf98c11c8e19c0b551021ee2cfa0408581195;
mem[373] = 144'hf8e003dfe94818abfdeb00d1f80917c1f683;
mem[374] = 144'hf9afee3902ca03d4e531044efdfa19b8fb91;
mem[375] = 144'hfec817caf228f1f313c4075f10e3f020e0c1;
mem[376] = 144'hf3d51cdce9d9f2241d5304c21b2ff502e7c1;
mem[377] = 144'he853e4d1068b14ff0be21814fb53e31bf677;
mem[378] = 144'hf4320efde68d0f6e00bde457f0b8066809c8;
mem[379] = 144'hf34f1a0df28805c9e9d301c813b20a010830;
mem[380] = 144'h1835e50ef67ce9f716801d38f75b0cbb0b7d;
mem[381] = 144'h0eb1fc78e8bceda7e418fb38fc040fcf0b9a;
mem[382] = 144'hf16ce3220072eef0feb5e7dffdddf1d9ffe3;
mem[383] = 144'h0eef14bf0ef01772ef000a130dbe1169f010;
mem[384] = 144'h070217c81e18f8b6fc67f579155d13400df5;
mem[385] = 144'he57fe8e0ef1aeb6c0323f8450afaf03de43b;
mem[386] = 144'h16431a39f5a60a7ff77ee2121f29fb32eba1;
mem[387] = 144'h049204e4e750eb34ef4003aa13bde1e8115e;
mem[388] = 144'h1c58fc2c0ee7eb7209c4f0611218effde594;
mem[389] = 144'h0ea0f37ee658ee830b8e1a7205b50f0bf7ea;
mem[390] = 144'h06370b5dfbf6fe38e0aff5cb1185e5ffff0e;
mem[391] = 144'he9db1012f37a166c1795f9e21e0ae4b0000c;
mem[392] = 144'hff71e73d0a79f36df47a0c781600e86c0b11;
mem[393] = 144'h14adf0781cd01b2c0280e552f4061cc9e1a1;
mem[394] = 144'h0d1ceacfee4bec251dbfe92c1a47e2271f51;
mem[395] = 144'hff1ef54cfd610cebe6fe16990689ed35016b;
mem[396] = 144'h1ff4e42afae3026ff76f0df6fe961244014f;
mem[397] = 144'hec3b0cfbf08b07171557e4130e531fda1f08;
mem[398] = 144'hf0ff1d77169417da10b1e919f22f10721850;
mem[399] = 144'hf71617630b3214ab0a091d3cf01ff8fcfc41;
mem[400] = 144'h09aafd0de01c001df58be013e4e612bbe32d;
mem[401] = 144'hf636f2531eeef3c71d2419ad13bf0e75106a;
mem[402] = 144'h004c05081e56024bef1e051ce11601611bc3;
mem[403] = 144'h0c2800f9fa0e10e81f03e2521f0f04a60298;
mem[404] = 144'hedb7085afe4218cc03530f0efbbae2c7f9a0;
mem[405] = 144'h10fd0ef9f3601e6111e60fec1faf0cf10ccf;
mem[406] = 144'h13970a5908c5f94b1f140b19f521f9700b6d;
mem[407] = 144'he781f94907c4ed86172bfe1c19f8f8e0fc62;
mem[408] = 144'h1fc704140d501909e85219b704fe01d0163f;
mem[409] = 144'h16c8e9ec02b213dc02fcfeb1f3d6ec5ff8dc;
mem[410] = 144'h02761c5110c5f6bb0306f968e4e61ba512e9;
mem[411] = 144'h139cfdd0e346e12fe34309dc1f191263177d;
mem[412] = 144'heac8e9b3eb59e50ee7841ba7f6540123fb5b;
mem[413] = 144'h037ffc32ee0a036218bf1bde0a45e95bf2aa;
mem[414] = 144'hfd7d1e05e2abf7f8fd07ff68e487fdb71381;
mem[415] = 144'hf13ffd36e17ee3841424e0e9fcdc009b09eb;
mem[416] = 144'hea8b14c3150de0d101bcee1a15d9eec5fbd7;
mem[417] = 144'he67ce4140d481a43e817f7f114a1ea670318;
mem[418] = 144'he08211a61d1b1510ebfd15e7e28c15c81c2c;
mem[419] = 144'h1951f6bd0b42fd66162f0ad7e98304a3f538;
mem[420] = 144'heae9f419f920ea3c1675f43204e2020305c4;
mem[421] = 144'hef67f5c51ef100a114f811e6e27416adfc41;
mem[422] = 144'h0ba4f36bee17e5661cd0f5b4ea600b64ed01;
mem[423] = 144'h0bc0eaa7053ce8a7ee5be078ec751d19168e;
mem[424] = 144'h1d28e87405481ea50f60ff59112beda5f20e;
mem[425] = 144'hffd5ec301de40e43fee6e7830e03ece8ec33;
mem[426] = 144'he868ef3ee387f20f037be458ffa81e66093d;
mem[427] = 144'h009c1a24e42be69b01f3fb67ecbdf19d0350;
mem[428] = 144'h1a720508f4291bb1fb69ef4af84f1bde0dde;
mem[429] = 144'hedc102a10276096e1ca2ebe6f16d0a661d02;
mem[430] = 144'hed06e805f167eed7ff93e083f6ec088f1390;
mem[431] = 144'h0f9eee1018a81681f807f8fce24ee26dfd18;
mem[432] = 144'h084decba0e91fc411e7b0d38f2effb3616dc;
mem[433] = 144'h07eb1f00f380ea86e518e4f4f08ef0311bdb;
mem[434] = 144'h1ad20a541f46f11c02ec03a4137a080005db;
mem[435] = 144'hf114173e02c106ca12d9165616980f780501;
mem[436] = 144'hf6331aff170ae643fb37fb0909a1eb47ec94;
mem[437] = 144'he23ee2c3e4f91494fb65f75df0f4e8911843;
mem[438] = 144'h1dae03ffe32bf1b0122df4ef052fe9c0f792;
mem[439] = 144'h16c102ad0c4f04050bfefbe8e9a0e189000e;
mem[440] = 144'h1422e70b066016871b67f0d416c819e810f5;
mem[441] = 144'h17c70953ea5ce921e6f90d760beef5a5fb0a;
mem[442] = 144'h10b71be7097bfa40ec67113de1dc00af1893;
mem[443] = 144'h14b6ece21e750907e956122f1701fff41f17;
mem[444] = 144'h1f1a0013e97ee9761aec08b0f3a10c45f5c0;
mem[445] = 144'h13f8fe3908f8fbeaf6a01ec5009de819fd60;
mem[446] = 144'h1f97f73d0ab414da0e38fe741decefeae4f3;
mem[447] = 144'h0ae5e4bd018817281ce51c5fecea055dec11;
mem[448] = 144'h1886145a1a42e105e60e1868e4e51c030da7;
mem[449] = 144'h1ef3e294ec13e27df79aee9f09daf5f20d52;
mem[450] = 144'hfa49fe0fea18eb46f05415c11707f055e00d;
mem[451] = 144'he463f604f6dbf74c199ee431ef45e4e716b0;
mem[452] = 144'h07b1ee4be3ad10bb04c30fe6e21d01670c99;
mem[453] = 144'h1cbefa18f0cded0800461da4f356e839ed05;
mem[454] = 144'hf2120972ed78f77ce4beedb1ef8de42d10a2;
mem[455] = 144'he935e148e92f0bf5f32cea26fdc305d5e72e;
mem[456] = 144'h1dc91360e17bffbff7820c11f937fb0dfe8a;
mem[457] = 144'h0d59126de0070e6c044003000369e17cf3d1;
mem[458] = 144'hfa57f5c9eac91448f140f9cc022be92fedc4;
mem[459] = 144'he5940c5e187117a4f738eeb3faa0e91310d5;
mem[460] = 144'h129eea56eb37ff9c0009073ce4680e70e673;
mem[461] = 144'h18db150903ed11e1fbebea351ebaef8afcbd;
mem[462] = 144'hf590f7061d36172c0a86fc40fc9c09ca086e;
mem[463] = 144'hf27dfb97f3dd066a0ac714af0343ee4507ca;
mem[464] = 144'h1bf2e030fe81e68be3a91d65f2950dccec78;
mem[465] = 144'h0971edabf9570453041f184317321d01e384;
mem[466] = 144'h0edfee11e030fb99f393ed1e043e19e719cb;
mem[467] = 144'hf413fd420a58f9b911edf717fab11262091d;
mem[468] = 144'hfbe3f7f8f89c1939112bf699f9db17c305f3;
mem[469] = 144'h01f0f49df72aec49088df692ed1bfd35e6c7;
mem[470] = 144'he0a90aa516f81305faa5f78be62be692e69c;
mem[471] = 144'hfc63e7b6f646f736111ffdca1a1718751294;
mem[472] = 144'hf5b519520ff11808e7ac1569e790ff0feaab;
mem[473] = 144'h0846e08117191162f6351c9e1832f74908a6;
mem[474] = 144'h109cefcc0100ed541b7dff8af794ea70fb2c;
mem[475] = 144'hee82f41a15cdeece163a1012f8fdfe7b0e76;
mem[476] = 144'h1473eb32f5ec1787e8880585fc2bec9a1ff7;
mem[477] = 144'h04cd188d1d8be7541184170aebb81c18ef57;
mem[478] = 144'h17dd10061e6ae364efb615220984fdf7e5e7;
mem[479] = 144'hf10c0efeea3aff9cf47e136be276f374fde3;
mem[480] = 144'heec90b6d094b0727f571e10d076de5f31f5c;
mem[481] = 144'h0e45fedd1242e5e4ec05ece104c7f8630f26;
mem[482] = 144'he9ac0691efe2fe71e0ff07c31043111b0bb4;
mem[483] = 144'h127eef390b6d0eba1589f084f4a1ec60fae3;
mem[484] = 144'hfa9df3b9e914efdb0287fc931d5f0745fdb5;
mem[485] = 144'he9e5f708092618f10e6e17e608a5f286ef0e;
mem[486] = 144'hf9fdffcce725e0bff6bffc11fa8de61f08de;
mem[487] = 144'he104088b07ec0beb14e513fbebeb05171bcd;
mem[488] = 144'h1836f27c0aba0d68ea1b1e35fc5ee5131113;
mem[489] = 144'h082e1ed7f46f0bdb149c0b3fe42bff3feaf7;
mem[490] = 144'hea490796f20be87fe697fbb7eb62e7521e13;
mem[491] = 144'h11490e1419d1fb91e8a6fb9ffc261df51b0e;
mem[492] = 144'h0403eae30e8cf3f4fd4418a003d2fbc00d3b;
mem[493] = 144'hfb9ae1a610d0f4b00f900925e8fbe8d71223;
mem[494] = 144'h1cce15e407aeff9918a70344f672fd73eb0e;
mem[495] = 144'h0ce7e116e82205a4e25a14f717da1fc3f651;
mem[496] = 144'h070814daf7d1eb6cf5661366e7e81bb90835;
mem[497] = 144'hf2f7f97eee8eedb4fb381b7d0877172ce1f9;
mem[498] = 144'h142debcbf62a12410599eb2301400403e4ba;
mem[499] = 144'hffe4115ae86b1d21f48dfbb0fbc701fa02f0;
mem[500] = 144'hf241e26ce2ec06391efee22c061df15fef6f;
mem[501] = 144'hf738e378e62b0ee1fa6d0f070dcc0aef0712;
mem[502] = 144'h16b8e2021dc1eeb31f22fddf14adf954105b;
mem[503] = 144'he5dcff0716f9f60e12ba02fe0acb0dd816c7;
mem[504] = 144'hf7de0432e08e1d03178117e9ee0b1d9e1d7d;
mem[505] = 144'h1afce080ec7e1c96fe73f1b9190beb4de6ba;
mem[506] = 144'h0a7c1b3309941595ebc00b8def8dfcf80a1f;
mem[507] = 144'he3aff7f3f7e81f34ed3010f60a20f08f17e5;
mem[508] = 144'h0ac1f81bf3f7e2481b12066a13911f810135;
mem[509] = 144'h0907f25fe3e41de810d2f397198fe5d415ba;
mem[510] = 144'he842f17f110d0d6f159f089b01cffa3bf272;
mem[511] = 144'hebce0298f952e5591093e4d401f71b820d19;
mem[512] = 144'h1e2d0d9cfb130dafffa9e7cf171df837178d;
mem[513] = 144'hfeb6fc900b15fd77ed4ffa7af3440512f11c;
mem[514] = 144'h1a37eca4eeefe85d1d9bf288057f196b1fc5;
mem[515] = 144'hfbf2f173fc22183e0f89f396f4f11b21ebaa;
mem[516] = 144'h19ed06bb0cace4e7e6c20e981bb816b1fa6b;
mem[517] = 144'hf19b0fade19a1024f6c8fb030232eebe0621;
mem[518] = 144'h1dca108ef9ed0bf31bf4f0e5ea271eed095b;
mem[519] = 144'h0b3a1f9dfe2a150c06fbe29efcc10dd1e9e9;
mem[520] = 144'heb6ae11c0984f089ff11f8cae787fe95ef35;
mem[521] = 144'h1ec813d01ff10db91eacfdbf07ee1522f369;
mem[522] = 144'he64f08c2f8c70b97ef8ee994046e02420642;
mem[523] = 144'h0b9b0f150e07eb48eda6ea04005bfd74ede4;
mem[524] = 144'h0703f3740207efe702b402ae00ddf75ce59b;
mem[525] = 144'hf67de4e106e41721032ae16cecf9e61cfd43;
mem[526] = 144'hfaa219a6f38904591dad158afc99106d0416;
mem[527] = 144'h0073e154e402f56f1cd916321f41f125e69b;
mem[528] = 144'h14d4f8e814141c5dfc1bf778fcc0ec0ee986;
mem[529] = 144'he05fe06cf96bed6bf901e7bff8a901e60e10;
mem[530] = 144'h11ca172b1060e3491664e12fec35f78ef420;
mem[531] = 144'heac701981bfa07060a871ddce6551f1bef1f;
mem[532] = 144'h0bb3157f1a77f10ff34407c51bf8ea141150;
mem[533] = 144'h0533e531f3f0f9d9f49100fbe4e1ed60023d;
mem[534] = 144'h1476126aebaae258e0f61929ed7c046f0ac6;
mem[535] = 144'h1c650a3b0c380a4ce937f207135af846e533;
mem[536] = 144'hf02bf379e9311b1fecd8e46be455eaf7e348;
mem[537] = 144'h0ae3e6f5ed76efb4e4050a7ae3ece198f43b;
mem[538] = 144'h11621eabfa4fefa60fa8077fe43d147cf3e5;
mem[539] = 144'h180ae41e1eef0dcfefc6f572e1060a310ad5;
mem[540] = 144'h1541fbbbf167f85116471799ec63f4f11a45;
mem[541] = 144'h1b8e1f2debd117be122f1ccee4bb12fcfaf6;
mem[542] = 144'hee21e26bf9c7164beb83efed0bc8e662efab;
mem[543] = 144'h0c81eb76f6f2194c0245ecc2000be982ec2a;
mem[544] = 144'h11a6e0bfe9000e0f18590f80105605200c7b;
mem[545] = 144'hfece0a4a097ee939fd6ffdccffec1f8ae8f3;
mem[546] = 144'h1075e80bee760829e0820ce50038f59d13ca;
mem[547] = 144'hf0ef01fe047f1df0f282e8510af51e6bed25;
mem[548] = 144'he6ac05a6f88c162af850e80d105ef09ae243;
mem[549] = 144'h0904f2ad1d120e32fd99f57ee9d1070409bb;
mem[550] = 144'hec14146404051254fe4ae339e625f1da05e7;
mem[551] = 144'hfda91e3be600f6be1afbe360070fe9df0835;
mem[552] = 144'h05271a2a09be105bf03205acffe7e3c2e70a;
mem[553] = 144'he96e1ad9f172ebd9ee1507c71ed30ab4e24a;
mem[554] = 144'he1711356e442091def9c0966ecea15fbe086;
mem[555] = 144'hf78b0a54e08ee1f0045c0e4109d4fae1e474;
mem[556] = 144'h19eb18b801601a2bf0affb73facf1851fde6;
mem[557] = 144'hefa2f5d7ffa5f16b15e304681240e8e2090d;
mem[558] = 144'hf437fdae0235e79ee42ef1a41f5f18a2144b;
mem[559] = 144'h1909e0d3fae0e2fc1d3de84be349e97ceafb;
mem[560] = 144'hf7f1ed41ef94ee0cf5b3e7e0098c081005b4;
mem[561] = 144'h1aa7f602e411ec8d1f1b103fedd2f9171e83;
mem[562] = 144'hf9ef0951fcb3e1dd08941cefe342079bfd88;
mem[563] = 144'h0bc517e604f80896f598edeae329f381f09f;
mem[564] = 144'he558f743ef8f0bc8fe41edca027e0aeb06e2;
mem[565] = 144'he79cfaaa19f1faae0a80e7560bc20731108e;
mem[566] = 144'he28df884fa670a4e197efcc2114e0acd0f62;
mem[567] = 144'h1d5c185ee3b0e539fb15f681fb1fea15e635;
mem[568] = 144'hfe0505fdf53e0a2e0d030aa3f84d13a81355;
mem[569] = 144'he224e1df1cb3f0b2047be62f194a0e94f0b0;
mem[570] = 144'hf26afee2f84be3fbfa551b5315b3f35d1f08;
mem[571] = 144'he1f1fce8fcf3ea0e1622f886fd6cf50ae5e6;
mem[572] = 144'h1412f7c01e2e169ce42be16afe661642031f;
mem[573] = 144'h1d27e9d6f00602600138f0831804e6930dc6;
mem[574] = 144'he06905ff1bbe133404bb14541dcb11bfe479;
mem[575] = 144'he094fbcdec7df0d208a1f1d4112ce88a18be;
mem[576] = 144'he094e97c1dc6e76ff268ffb7ed85fb91e9de;
mem[577] = 144'h0e74eccbf98fe011e49d07b2f68e0de20eb4;
mem[578] = 144'h0cecfbfdf09be8b7f6ff0ff0e397e5900594;
mem[579] = 144'h14441c0210ef11bf1a27192decdd103c1c54;
mem[580] = 144'he0dbe8f41a0eff32ee3ff3bc14c1ee76e516;
mem[581] = 144'he1f70cca0e9e1f240958125af55d1faff394;
mem[582] = 144'h0679f6a312761054e935192c1ef007a7fdb4;
mem[583] = 144'hffe80d1714d00671e83ae8f8fd9bfd9be224;
mem[584] = 144'h0ec0053a0951ee5e1117f136ea9ee0bff8f4;
mem[585] = 144'hedb306e0e0fee507f2d60f6df366e3aff552;
mem[586] = 144'h0d2d058b01cc0dabf0f1e4380e561787edfb;
mem[587] = 144'hf5ca0190f2d20a21039de506f13215b61bd7;
mem[588] = 144'h17cce4dbe3e60e4706c5faebf5f7069ce240;
mem[589] = 144'hfc4b0d60fbae0174fe89eaad028dfe8d141e;
mem[590] = 144'h05c509dced09f810fbdaeac5f3b7f83c19e8;
mem[591] = 144'hf85ce41bf31f0cba059df344f088e5aae728;
mem[592] = 144'h09a906cbf293f18b12bfedc6f3d01145024a;
mem[593] = 144'h029815eb191009e6104a07fa0b4de54a0f7e;
mem[594] = 144'h04310735f6220c74e74d106ef574f809fe91;
mem[595] = 144'h0d2de328efd31981e21007cafff6ed3b0910;
mem[596] = 144'h1acde7750ceef6d6f487e1fbe0b014ddfa96;
mem[597] = 144'hfecaeed20a1c0282f630febd16171f61f2d5;
mem[598] = 144'h0e92f604e5020125f00a1a91fcb91ad8e92a;
mem[599] = 144'h120fe55de5e8198ae4f9f75b1c53e259f4b3;
mem[600] = 144'h14a617a3072b147aff6a08d5139decca0497;
mem[601] = 144'hf58a0e7018c7e218f6ac16ee02e106e01de7;
mem[602] = 144'h13ff13d3fd041fd6fe1a1cb010c400670ee1;
mem[603] = 144'h02eb14ea074206eeefdfe3291da201cc0757;
mem[604] = 144'h1d670b5df003e7c8f4c203bffd0afd52e7da;
mem[605] = 144'h00fef22f006bee07fc86fc7f0351e55be205;
mem[606] = 144'h00c8093a079f1f73e4961e55ecc7f7c60edc;
mem[607] = 144'hf4480d510b48f49a02fc18adeeec0e2a0166;
mem[608] = 144'hf2ea1abceb74012414ec0e6cfcaee766ec66;
mem[609] = 144'h1b0c1a8817bb108af5ae18991b16e4aa026f;
mem[610] = 144'h056c0f3319ca0101029d02b10861ebfe035b;
mem[611] = 144'h04e71ea30c66ee800c91f97bf1a0171f150f;
mem[612] = 144'hf7861ecc1952eda7ee85ece50fc7f4be1f12;
mem[613] = 144'hea1012ec073efb1c056ee8ce1c7e0e2a012f;
mem[614] = 144'he39c0c1de15f1f5fe7e8ea02e800ecbbf464;
mem[615] = 144'h0af4fc4ded321cf4041cec901a140e2d0941;
mem[616] = 144'h12d4154d13befbb81ab31137dfd60d43e95f;
mem[617] = 144'h03c1e49d09d7fee7ffd70b1ef62ae08bfb7e;
mem[618] = 144'h0e1df8a105c80d98f897e319f4ad04ae134a;
mem[619] = 144'hfb951ec8fc630a22ecebeea7e0651da40d0b;
mem[620] = 144'hf8bf1d0aedddfd70ee860e63e4f4ecdefce7;
mem[621] = 144'h104a05cbe376f78f0d59eb4e0cb005d60032;
mem[622] = 144'h0672feb00d97180509aff097163efb9beccb;
mem[623] = 144'h128706950a2005fde946070fe6d1171fffd2;
mem[624] = 144'hef5a09cce1231c90ea300c3d0ee31c7b0f69;
mem[625] = 144'h1dc50029f9a8f65115a31d091ca1f9641289;
mem[626] = 144'hf613f369e0d002bafaa7f20d191613e0eb39;
mem[627] = 144'h1fa4087df2e0e67bed5df6cafade0a1bf8e2;
mem[628] = 144'hfb0202ab1caceea5e165e451e698ff4215ee;
mem[629] = 144'h1bdb10c6ed9ee48d1636fef00ff914f80e1a;
mem[630] = 144'h13c7f8c515ceeb670d240591efa4e30a1647;
mem[631] = 144'hf846e04312c8fb9ae8eaf2c706dd10210569;
mem[632] = 144'hf743e98318b9f8f807b0093100cd001f0065;
mem[633] = 144'hf9ec0e6b1d1efa1619940d1df74c09ac0ea3;
mem[634] = 144'h14c30a2d1de61d70ed5deae90e07e892066f;
mem[635] = 144'h1027ffaa1866fccf058d114fea031e501d97;
mem[636] = 144'h070bff4cf1e0f93af916096f13111b7deb55;
mem[637] = 144'hecd0ef85eb8509a31019e468173ce97a1856;
mem[638] = 144'h187a0434e311171d0d2de69a030c111e0acf;
mem[639] = 144'he7ce135f0eea1260fb0319c7fb4d041715a2;
mem[640] = 144'h1ca0f09c106feaa1e0f6ff801801e58bf2a0;
mem[641] = 144'he2ab0106f6c3f9eaf9561159fac9f7401a28;
mem[642] = 144'h0d12e2c0e87613be0118efac0b190e490595;
mem[643] = 144'hfd82e4a10483150214bf09610633e687eac7;
mem[644] = 144'h04d8e5891bf310f2e0fde002e31910e1e35b;
mem[645] = 144'hfa42f5aa0d381620eb5f19e6e197f7691a54;
mem[646] = 144'hf95ae13de7aefbf8f524fc70171d0ceb0a2c;
mem[647] = 144'he4610b690b8e1afde7b30fda17fafcb80b06;
mem[648] = 144'he944e3420e41fe85ee51092cf1d314a51c85;
mem[649] = 144'he2fd1a65f87efdfbff48e5ef00bbfc3eec42;
mem[650] = 144'h18e1070be602123ee4f40203ed9a1b5ce988;
mem[651] = 144'hf1ce0761f814ec9d024b124b0212e6ff13ea;
mem[652] = 144'hed4ce86714d906950a47f26ded9ce0fcf8c6;
mem[653] = 144'h188d1bc8fc2df1d4139ff7f6177d19fdfd2a;
mem[654] = 144'h088b126605c61edb06effd12181311d4024e;
mem[655] = 144'he8e7f48804f6161d0931099ef7c4fb62020f;
mem[656] = 144'h18871844f0b11e52fd2bfefae73ceb2f1d53;
mem[657] = 144'h0f940597112bf4cae7920afe1fb211af1e7e;
mem[658] = 144'hea4c1579f8d612cc18b6f2530bdb0b2ee9e8;
mem[659] = 144'hff93ed8e08a1fb2bedf80eebe32505270f5e;
mem[660] = 144'hebe8f0641fcbf95a122b08bbebe20f360e90;
mem[661] = 144'hf9e1eea3ebfc0a14f2f6fc1a0f9ce94bf4b8;
mem[662] = 144'he3befcd51cb4085ce6711e38e415ea07f8e3;
mem[663] = 144'h09501182fe0d03d7f8261266f49af24212b6;
mem[664] = 144'he9cd18050378f1411470f276f379ea9b19ac;
mem[665] = 144'hfffa0c8c0661082de378f8b11345070aef1b;
mem[666] = 144'hf5ff0302e3baeff11c37e90cf2e3e074ea92;
mem[667] = 144'h1d40f9000dd3ed42e8e8097c166208ca0ba8;
mem[668] = 144'h0535120af57d1c18e2ddf0a4ea0cebc3ed48;
mem[669] = 144'hf9cde970f70211271b69fcb2efb3f6561eab;
mem[670] = 144'h1a95156106d4e5c70635f1fd1eebfd95e964;
mem[671] = 144'h196b1b070531f40ae670f34f036a131dee5f;
mem[672] = 144'h0c7c0b00ff33edae18fa02e01302f8fd1402;
mem[673] = 144'h14b2fa371186fe1fe1181db21849174307f0;
mem[674] = 144'he019f7a315cd001fe9901da40c871a7ffc82;
mem[675] = 144'hf189f708f9870e89e6610ed418bf1daa17dc;
mem[676] = 144'he16ced6df96814a6e1321360fe4308b5e75b;
mem[677] = 144'he9ce0d5d1934f782e2ef0a15f58d1214ee67;
mem[678] = 144'h07c3f1e2072e0b1dee2a11bce3e10af31ab0;
mem[679] = 144'hfc601a5c19751bde1fb21fa01169e91cf855;
mem[680] = 144'hf721fade0c7605afeadc127609b11614fab3;
mem[681] = 144'hfc7418c7f030f2bceb4de378fe81e9ca0589;
mem[682] = 144'hfe42ecf61785e072016af05cf43becd0f66b;
mem[683] = 144'h1a7bfbb6fe47f64ce2f40fe2ead415e2f667;
mem[684] = 144'hebbff640ee2e0410015f0a41f74d1f55f677;
mem[685] = 144'he3e6ffc70dc7e938fd8ef5b0ee6ef3130e41;
mem[686] = 144'hf2d10e39eba7fb610dd1faa2e23b0c1efb66;
mem[687] = 144'h0b59ee2e077d1b5ffa0cfbbbe8860b89e1a0;
mem[688] = 144'he0c2fa0a1d4c06c5f3b0e363e4160a1eee4c;
mem[689] = 144'he795148c0245e82ef56de6810013ed540b9f;
mem[690] = 144'h03f80a53eda6f1b4fbd2eec41330148a0268;
mem[691] = 144'h09e9fb47efec1bf407a61d5216ec1610f6c1;
mem[692] = 144'h0a1df4230a3c019a19c6f93de09eeff2ff10;
mem[693] = 144'h17cff9e0e3ab0cc61324fd64133f0953e76e;
mem[694] = 144'hea17f4cef0be1ab616271cfbf09ae40f01bc;
mem[695] = 144'he941f69bfa24dffaf62517cef63eff64e50c;
mem[696] = 144'hff49e94303201e0e1acef26efd16f2f9fd14;
mem[697] = 144'hf392065d0668e6b0fa0c12711f52e94408e5;
mem[698] = 144'h0b1101f50c8602c7f1ef1905ec69eb1f0cff;
mem[699] = 144'h1ca9f496f1740d0bfee50d03e56113fe125f;
mem[700] = 144'h0c97f7eeeaa106dae223e03f03bd12c01753;
mem[701] = 144'h0595106f14ed04e71e44facfe773fceb0ce5;
mem[702] = 144'h0a60edeaff02013ef459e0d3f81d1b4f1ba1;
mem[703] = 144'hf708ea8df11e05d813800558edcdeda40220;
mem[704] = 144'hfeec06150245e96a1f7715cbf8b703f2ed0b;
mem[705] = 144'h075f0b6ee4a9ebe603140d760692fa4df4ac;
mem[706] = 144'h02fa19531bdbe7a9e3c702630a47031efd90;
mem[707] = 144'hfa0d10811bdcf2fae6a5e2f1e5711032eb72;
mem[708] = 144'hfd5b19d714abe693ec95f0d116ec0eff1797;
mem[709] = 144'h18091c50f4a4f18212f1e758ea961f71f4bf;
mem[710] = 144'hf49de2b30c821a161269eef4fc42e1c7ea2b;
mem[711] = 144'he4a102c70a1ffbac1a12ed14f3bef742fbca;
mem[712] = 144'hff7fee40fa11185d119e1d4907b10537f48d;
mem[713] = 144'h16da1e59ed0002180990ebc4f7ce1e74fb63;
mem[714] = 144'he70d051d16281fd7faaf0e11f1451e50e041;
mem[715] = 144'h08380a4b0bbce6740b97f5ebed8efe5402d6;
mem[716] = 144'h0e99eb51f3f20b98e2b4e92df3b8ed590c27;
mem[717] = 144'hf2e61cb215741c210485ea42ea140bdef7ad;
mem[718] = 144'h0700e4d7f0250580f495ff8affa4fa95ec14;
mem[719] = 144'h1277f90c083201e70bf219841a5cf74e08bd;
mem[720] = 144'hf8c1f425e6f71638e9c3f641f4b0fad41c1e;
mem[721] = 144'he6fe17f3f0111ad210d8f44de1540223fd1b;
mem[722] = 144'h0341f18b1e1118bef863ed1f0147e0ff1562;
mem[723] = 144'hf3351aa4fcc2f3fb1324fb29eb5e0d021fc6;
mem[724] = 144'heccd015307d5e31906fbf22afe4ef5bae112;
mem[725] = 144'he6240a1616c8e947f95ff66808cc1198e29b;
mem[726] = 144'hf14d039f01ede418ec00e4400b7b16090c5a;
mem[727] = 144'h11370a071d8306c4fe34edbc142c122c1249;
mem[728] = 144'hfba3f3feeabc1dae1af6fb0ef91f1e59e664;
mem[729] = 144'h02df14120bcb1a92ff63f60516450ebb090e;
mem[730] = 144'he8caeeee066307c8f0eff985e3f90759e9c6;
mem[731] = 144'hed430a72f50204c7e4b513ebed53ef5fef40;
mem[732] = 144'h0416e869f6e1f025007e0ebcfdf216340d95;
mem[733] = 144'h0795efce111ce4d4f688e9f019e6e264116f;
mem[734] = 144'hf99b09ffe4caf206ee961aaa14c81051ed52;
mem[735] = 144'hef42fdac09d4ee131557e8e811591554febf;
mem[736] = 144'hf58b03290c6bf4aded1ff3790e9ce52ae342;
mem[737] = 144'h0af31b990a5718050f9308df174fe5cd130c;
mem[738] = 144'h0c731fdef8041e190e3bfbc7f53be60f1fc1;
mem[739] = 144'h06bf084d0209032e19cae094e0dcefc81d62;
mem[740] = 144'hec94ea620cd51c1701770dace999f3611469;
mem[741] = 144'hf54de69ce7c5f381f479f30fe92a1e1af51b;
mem[742] = 144'h02a8f807083e08c8f93eee9cf0b710191220;
mem[743] = 144'heb59eb5cf3511291f0df1c4e0194e8e8f382;
mem[744] = 144'he58610d8eea600f6ee6afc9af1ca16fcfb95;
mem[745] = 144'hf6ac1deae9b507201bf7e523e22be14e18e3;
mem[746] = 144'h15b21fea1271f0fa0193e298faebff0f1cfb;
mem[747] = 144'h16f4011f179715731cf3ef6ef955e739e3e6;
mem[748] = 144'he450fd24f4bb02530d0b05ee01651bcce1fe;
mem[749] = 144'h0cfb0bf516a6033de86f1a4ceced0afde61f;
mem[750] = 144'hea610cb205d8f1221acbe0220477e1690552;
mem[751] = 144'hf81900bd166bf04fe1461218fc4d1a17077e;
mem[752] = 144'he2bd1cbef471062e1b971e8fe68e0de71414;
mem[753] = 144'h01c1146bfe4a07b1fad4ed90e9e6174a1225;
mem[754] = 144'h1b5c15661f081c52e616e91a1bc900f21e39;
mem[755] = 144'h12a31d2e08a1035df4000d0b05c2e28ee9fc;
mem[756] = 144'h0c64e931ff5407580d3bec6defb6e823122b;
mem[757] = 144'h0c6211f91001e72a1f7be053147de956e6f4;
mem[758] = 144'h16a51fe607b9fecaf09e12030c8ee642162c;
mem[759] = 144'hedc71f070e641e4bf0460aaff7450fc50efa;
mem[760] = 144'h1119f411e7eb00a2fbfcf6bde9630e29f426;
mem[761] = 144'he57efc36f5241889198f146511b4f49f09ea;
mem[762] = 144'hf936f427f71206d8f9f91e61164102fe1f85;
mem[763] = 144'h0e57fcfe0effe3b1f1e402ea01f5ed9d0c34;
mem[764] = 144'he3731a09f1cbe917fee9eeebe363e6e2057d;
mem[765] = 144'h1b66e10c14db17460169edde0ae80edee941;
mem[766] = 144'h024f0147150810f5161216450b88167af1cd;
mem[767] = 144'h13481c99e070038bedb1e2e911bd0b1a09ce;
mem[768] = 144'h1b98fbdbf811fb3f0118f73d1ec11930e0c1;
mem[769] = 144'h15a619cd186fff3efc95fd11105ceb7f05a9;
mem[770] = 144'h1c6e12a5e7d008d70ab3f80aefc61cf50fbd;
mem[771] = 144'h1e2310540ac208fcf20611fa0d4efd931b74;
mem[772] = 144'h0fd6e41900901f7bf69b0520e3a2e0a6ec66;
mem[773] = 144'heaf00ca3fe401eed0342eaa9eb6c0df50571;
mem[774] = 144'hfba901e50e16f26706521dc0038eed58fd44;
mem[775] = 144'h04afe02d101f1633ea37e5bf08e707b8e66a;
mem[776] = 144'h0069e14decc6038f09e4f1ae01150b011f38;
mem[777] = 144'hfa060ccd1188f4a90a3fea4bf548f7abf859;
mem[778] = 144'h1525ecf819731bca036e0bcff67a0cacf71d;
mem[779] = 144'he240fd8a05b2e4580ca5f9cde39911011b28;
mem[780] = 144'hfe3bf896f2ea07e70f07fb96e73ae9b7037c;
mem[781] = 144'he39e1a8716e9f053e50b19c91513e74be606;
mem[782] = 144'h1b2e1672f2e814c3ff6410d41959e7a711e1;
mem[783] = 144'he0511d5f0a54ffdcffe8f60a171a1f380330;
mem[784] = 144'hff9804f5ee2bfd07e7e1062915741161e57d;
mem[785] = 144'hecedf4d10e02099d04cd002f1f3ce5681363;
mem[786] = 144'h19cf0a0610b4e5ccf2f812ca00b815f5eccc;
mem[787] = 144'h117f01acfc19062fe06f04261092e783fb2c;
mem[788] = 144'h02c616b311e7fe841092efd7ed231b321a6c;
mem[789] = 144'hf624e6e6f35d13e4e0ef17f9eb7bf26618b6;
mem[790] = 144'h04ff18bee2e40e2e0abeee62e2c1e591e5b2;
mem[791] = 144'h08bcec88ebe11fdb03d8ff4cec6b1a19eb0f;
mem[792] = 144'h1b7a1520e3fc16611fe51cf601351323fbc7;
mem[793] = 144'hfdb806fdf5ecee53153611f4f0a8ecfef375;
mem[794] = 144'he161f0c4e82903b1f153fc731b39e832f50e;
mem[795] = 144'hfa12fef60bcce75ce8eb01d012bef5efe976;
mem[796] = 144'hf2041ca5f87302161be0fc5bebed02cb1d7a;
mem[797] = 144'h0adc19e0ed5af1fc04e11a1ff2b9fac906a2;
mem[798] = 144'h10c31b64eee3160af0a70772f7e1e8b2eef7;
mem[799] = 144'hf197fdc41de5e5fd011a0facf825fdec0734;
mem[800] = 144'hf120095cf94518d8f775fbc01265059b0dd9;
mem[801] = 144'hf929eae61cecf757e1db0e230c91e7df184c;
mem[802] = 144'h06aa02cc0514e4c8064f14050f611bd7e253;
mem[803] = 144'h06661668eb12ea51ffbce17eedb2ea58ee47;
mem[804] = 144'h01a81e5de2971ee4005b1be6fdcb1a3e0bc2;
mem[805] = 144'hf747ed22068cfdf016fd0f0be9b006981982;
mem[806] = 144'he83913d4138a0050e4e41896ea671751e8ae;
mem[807] = 144'hee0dfdf70460096dec67e9d80ea00de81b35;
mem[808] = 144'h03441f6d190315b9e348f421031c1374f9b0;
mem[809] = 144'hee1ff913e40c0eb517381e0c098aff77f2fd;
mem[810] = 144'h1e5f143e04d4f60312b513f90ac9f6fa0790;
mem[811] = 144'h07391d381722e2af1bdd1ddaffc5ea790e87;
mem[812] = 144'h16301d00173ae45b1cb01140072e16841ac7;
mem[813] = 144'hfd50f4e616f20b631e6bfe6018880b91efd2;
mem[814] = 144'h11d7e4cde357e7420e79e0580d09f4dee8ab;
mem[815] = 144'h19d10053fd37fa54140c1773ebc809e80557;
mem[816] = 144'h0c70f9451982e0d1f1480c37fe1deeb11ee6;
mem[817] = 144'h0ba6ed901edc1306e0750290e416080213e3;
mem[818] = 144'h1b47f8bf07c1ebade9b819d8f0441e4cec12;
mem[819] = 144'hfcbe143a0c71fabf1f43e07c1dd6fadde8bb;
mem[820] = 144'hfa081b7519aa049d11020422fd81f87518db;
mem[821] = 144'hf5de1bbeed98f8590601e479fbd1fdf60244;
mem[822] = 144'h0538f4c8f93f0b59f9221c99058ce1930490;
mem[823] = 144'hfc9503a4e3e9ea04e64d1809f0d3e7861276;
mem[824] = 144'hee581eac0ec2e838f261f084fdfcf666f944;
mem[825] = 144'he473e8830eadf682f6a2f8131dd7e9a818bb;
mem[826] = 144'he6cb18250e25fbebe20a1a45042bf2370094;
mem[827] = 144'hfc8f1fb0e33ef2500e64ff2ff77cfce1fd73;
mem[828] = 144'h0a131f2b0d10e1d7075c1f191f17fdd0108d;
mem[829] = 144'h1da017d5e1f8ea861c9efa2f07bafcc40f93;
mem[830] = 144'h117af7fde6a60df71486e1f8108b187a1153;
mem[831] = 144'h19591594efe00ab2173e1fab07691411150f;
mem[832] = 144'hfa8e17921b1dfb7a13ef0289e0f808880527;
mem[833] = 144'h1b510c9aec13199bfe17e9dd06c4060e1f85;
mem[834] = 144'he77c149fff5be207fbee0296161ef7d704f7;
mem[835] = 144'he9d3e8751b32f79f0f3a1f4bff000aa2f0a7;
mem[836] = 144'h03a5fa360edaeee1f734184cf6780ce40da0;
mem[837] = 144'h1a98ed1a0c880c511721e98d185204651055;
mem[838] = 144'h0b21f107ea90135aeed2ec00009df01a07e8;
mem[839] = 144'h0d63f0430bbbe1c7f33818a1ef3d17b911d8;
mem[840] = 144'h0bfa06bee7cff02eea3ae315090ae165ea69;
mem[841] = 144'h0e46098e0644f807f95413700563160be9a0;
mem[842] = 144'h0dd008ee0dff0f450b8fed07eaef18bb045c;
mem[843] = 144'h0897f0d0e302eeda0fdce6be07c2f16cf135;
mem[844] = 144'h1dccffd90faeec271be10e2a17170044ef44;
mem[845] = 144'he594057ee2f1f558e67f1ebdfea4f6bdf58c;
mem[846] = 144'hf54eeb43103112931f49f012ef6600b6e01e;
mem[847] = 144'he62bebefe8c6ef39e591f0c4144a05a50155;
mem[848] = 144'h1a0a0e5f04e31b95049705dced37e529e342;
mem[849] = 144'hf7d604b1eb870bf1e6cbe7ce1f3518e604b6;
mem[850] = 144'hf5d0061aee1c0e65e0d014580271f48a0836;
mem[851] = 144'hed8510b0f7b8e523f3e3ece8e3ff1e4802d8;
mem[852] = 144'h0ec319b40769e77d1b331f88fc390b08ff08;
mem[853] = 144'heaf5e298f2f2e6b511bb1c23fff81a95faab;
mem[854] = 144'h1581f1ac196d0bbc1c8e07bd1ff507600c9e;
mem[855] = 144'he1291fad0acc1ca2eece0a31016ee4391826;
mem[856] = 144'hf200050fec67f57f1ae9f2e2f8840399fab8;
mem[857] = 144'heda803b4e2bdf2b4e3f0e98d177a01e919eb;
mem[858] = 144'h1d371a500d83ef0117d8055eff5cea561a08;
mem[859] = 144'hf03411c819b31ab7fa48fbb8fc19008311e7;
mem[860] = 144'h0e1ce1e4ef47ed72ff3715ccf3731fc80d2e;
mem[861] = 144'h13750a8c026cef0afb0c0df8082105ab10a9;
mem[862] = 144'he462e7880e68fcd4065d16ed00db05d31913;
mem[863] = 144'he5c1f0a303a8ed230e280f53fb8ce3950a63;
mem[864] = 144'heff1e0c3e411f906fafc12b2f303f02509b0;
mem[865] = 144'h1869e358f70d07091dca023bf43cfe2effea;
mem[866] = 144'he25a1206e93ae93aeea80d571a401221f758;
mem[867] = 144'h0cd3078108e2ef20066d14b2eb6cf1e6e543;
mem[868] = 144'hf2c9ff021055e85819ac1c8ff515e82c1553;
mem[869] = 144'hec79031cec7de1d1e6e718ce04b6fabde18b;
mem[870] = 144'h08cd114b1982e764f75b17b91f4cfe6bfa9b;
mem[871] = 144'h03aefcc4e8d9e6d8072ae2491450e07a1a5e;
mem[872] = 144'h1756f733f96f0ec6e786e7b9ed79ef680090;
mem[873] = 144'hf354f36112d5f59b055918c101b6064c0103;
mem[874] = 144'h158104261281eb5b1f791d461c7ffa4e0a4d;
mem[875] = 144'he9ab1b8ee499f7faf1a01b770ce719d5034a;
mem[876] = 144'hf46f16a7e815fbcc0387e7aeebfbec22eaa1;
mem[877] = 144'hee2b0bfcff5311a40adaefabfffafcd61535;
mem[878] = 144'h1b11072bfbd8e7401125fc25f0b91e97e5ee;
mem[879] = 144'he756060ef4870ad6188bed7c00a2e3a30e75;
mem[880] = 144'hf4cdfda5ee9e0d2011f00de60ac708aef532;
mem[881] = 144'hea07ee8905c60f211bcbffc8ef6f09d5e22c;
mem[882] = 144'h02751f3608a708b3f0e0e2c4f672ed9508bd;
mem[883] = 144'h1d32f97318f11fa31207f71af5a602020648;
mem[884] = 144'h1236fe0ff2350f7a034ffe9e049decdde5cf;
mem[885] = 144'h1dc3e03af4a1ecbff93bf4bae590e5adecd0;
mem[886] = 144'hed2d1e6915cf1d4af28cf38e10ca0f2ce8dc;
mem[887] = 144'h02fde373192403eafe831d2dfafdf3901b89;
mem[888] = 144'hf1ad17bb0e700b98e4940f98e269f73ff20e;
mem[889] = 144'h04d0e3171302156c0ef9ffaefa5cf410f590;
mem[890] = 144'hf9790493ff71ea1012fef1950b8f0ce31251;
mem[891] = 144'he036ece3f7f007f7f1ea1c68e398fc610b66;
mem[892] = 144'h1e65e029f375004bf2faec461a6bf1a0f73b;
mem[893] = 144'hf0190be2f6f5fba713b4ecdb11cb0cf90ffa;
mem[894] = 144'he2f10e5fe79d129ae9bd113de15e0262e09f;
mem[895] = 144'h1e2bfe50176714bc1771033b0e691e85e631;
mem[896] = 144'hf35107260624f6ae1333e4d31141f104ec8f;
mem[897] = 144'h03a617861b2e1127020bf2d1ec1301a8133b;
mem[898] = 144'h0f2f1273135b128d00bbe9571bdc1d63190b;
mem[899] = 144'h08ab15d6fee81a32e723fd85185a1b90e1de;
mem[900] = 144'he4daeabeed33e8da0158e8001f8319c8e1a2;
mem[901] = 144'hfd7c04d91bbbf0dd1e74fda0fc66111dee80;
mem[902] = 144'h19ba08fd0634f577e610ead9eee7ec71f3d8;
mem[903] = 144'he09d0c91eadc10fa1b70094a081af95af9db;
mem[904] = 144'h090114b3f7eef4ee0935f0c91979fb0409bb;
mem[905] = 144'h10b30d481ae71b931a46e9f4028df5ede32a;
mem[906] = 144'h12060f25f7830e9609a4f6b6178df906f159;
mem[907] = 144'he08b1f9be742ff64154be4d2ec4914dd0ee3;
mem[908] = 144'h0304106a1564e12915bc0f7cf0bef819e5a5;
mem[909] = 144'he7deff1cf41af85817100c3e1dbae018f4a5;
mem[910] = 144'hf031027ff99d1d5a0c13f76617b0fdfc12c2;
mem[911] = 144'h002d152a0de4e68901e0e74ae92f1377e1ca;
mem[912] = 144'h1830e7b50e241f260efa0441fa5d1d84e6e3;
mem[913] = 144'h1ce5f6c7e02d11f2ee7015b8fd6a111d189e;
mem[914] = 144'heb9916960adb043dedc4eeef1b5f1b88f039;
mem[915] = 144'h18f3e26d0849129c0514e709e2b7eaa4fd1d;
mem[916] = 144'hfe30e54e09bdebfaeb75e41b0df11914f57d;
mem[917] = 144'h0e87fc6a0aa21f3000590d5f0cc2f7c203b8;
mem[918] = 144'hf8f715e2fa8ef45c08d60d100e6b02d60d95;
mem[919] = 144'hfcf4ef2e02b4026ffb2ce51feb06f20ef272;
mem[920] = 144'h0103f17df221f70dfd4514fbe2c3086807c7;
mem[921] = 144'h1429e7ca03f00a17ff620b00f21bfd5515bd;
mem[922] = 144'hfe22e74f12490b44023d1c201e52154eebaa;
mem[923] = 144'hf527124b0c490d82ecdd12801959e157f58f;
mem[924] = 144'h026df0d1fe180c64006ff9c20ae4e2b9edb1;
mem[925] = 144'hf912f092f9070923105be4fc13d201fe138f;
mem[926] = 144'hf2a20ebaff69117e14d50c940a1efbaafdb9;
mem[927] = 144'h1ac8e382e10ce03318261f8afff407a60016;
mem[928] = 144'hf943e1281a86e778f456001bed770dad0237;
mem[929] = 144'he2570c761b3117ef0face706edafe5ac03da;
mem[930] = 144'hfb48ff14fe2ff828f627efca059df768f253;
mem[931] = 144'hedd7e624fdc0e8a617b41200f6bf1282f547;
mem[932] = 144'hf98c08861b66f96006f9f8bff71bf82cff2a;
mem[933] = 144'he59116261008ed39f919fb411ebeff39e4ef;
mem[934] = 144'h1908163603a90ac5ff76055a0aaafd1bed8d;
mem[935] = 144'hf57bf327e242fe2606f5f1fe0a0d097a112e;
mem[936] = 144'h0db5fe5ae6c3f51df9781080f2a716190d59;
mem[937] = 144'hff201970e8b91333f5ca07530b7ee4341ad6;
mem[938] = 144'hf4e2f663e59ce313f26403b2fbac16f11593;
mem[939] = 144'hfa8001d61b391cf3f8a809e903d0e2f8e867;
mem[940] = 144'h14951876ed0de941f939fb16f1c2e786ef69;
mem[941] = 144'h1360ecabeeeb0dba15b5189bfbc9027afb6e;
mem[942] = 144'he35e1e8aff8fe66310ddeedd18c8ede3ffff;
mem[943] = 144'hf71af8a1086ae613f2ff1386eebef115f969;
mem[944] = 144'he920e568fd89f401f956ffbee3a3f6a4e05b;
mem[945] = 144'hfa7c0194eb3efac61843ea42f394ef6bece7;
mem[946] = 144'he64817ec1c7214950fdceae6e683f613e807;
mem[947] = 144'h0bbf1ca5e6fc03390c25fd050901e6951c65;
mem[948] = 144'h1a50f3e7137ef5810e9703ba04a8f003ee6c;
mem[949] = 144'hedcc05b21e32e36d0388023bf6d7f2aafade;
mem[950] = 144'h04730331028be965f0f4fd0a07751de10ef5;
mem[951] = 144'hf617f04c14180d49e4c010edf2d6f0891c67;
mem[952] = 144'hff22e41512e9fdd813c0f030e3d317a9f030;
mem[953] = 144'hfdfbe362f578f28af03a06bef9f7f2d11c36;
mem[954] = 144'hef41ff23fad70ca3e64c085c124e0ca7e326;
mem[955] = 144'h16c70a89f207ec391c1e1a37ef2b09cee561;
mem[956] = 144'hfb6ffd3903e41f290a2eff41e898ff7eefaf;
mem[957] = 144'he137feda09561ab81043f7cdf22a0f7800a9;
mem[958] = 144'h14b8f157f48ce450e1e1f1ce1be90b9ce1d9;
mem[959] = 144'he15be6c5f99cf0d81057ff79ec6fe066ff2c;
mem[960] = 144'heb0a051dea9d115ff7e0176af529f1eae45f;
mem[961] = 144'h0193f340e209f900ee430130fa3efe06028c;
mem[962] = 144'hf368f55e05dbf383fa79ef0bf77b0c5501d4;
mem[963] = 144'hf42af958e73de372ef8df30414fc188df366;
mem[964] = 144'hfb65fdd9f66efd5c180f1b09f85706930380;
mem[965] = 144'h0484e368fb62e5831e6d1cd0e760072d04f8;
mem[966] = 144'he106f0250df0f1cb0ee6fd0616b7f4b8f8e9;
mem[967] = 144'hfbebe5940616f19ee19bec891f4d1f1af1e1;
mem[968] = 144'hee70e0b400bd17c0e3e70c47e6071cacff61;
mem[969] = 144'h0007f0e304c31eba17031158e89f0c1df35a;
mem[970] = 144'heac5e7461ff6e13805c114b10644f417e861;
mem[971] = 144'h07a2e80204a905b41f0b1866038316441250;
mem[972] = 144'h1fa7f66d10451d61e35e16d6e535f39d0743;
mem[973] = 144'h13891f6be9d3f3c3044a09cf12e918e7e92a;
mem[974] = 144'hfc010cddeacbf02ceea0108afbc81b3d125a;
mem[975] = 144'h15a31cb9f0d9f7b51a6a0521fb4ee69ffded;
mem[976] = 144'he56913edf6131a68fa8fe16c1762e0b0f1be;
mem[977] = 144'he9ecfc5cfd4f17acfacbe9d7f82cfe460235;
mem[978] = 144'h11eeed24ee83f471e391f1a1f1a70ddd1487;
mem[979] = 144'he1a00211e6e80b4df5eff6f0e2db016cfb68;
mem[980] = 144'h1c7ced82f14be696fe4b1bccf7d008070b98;
mem[981] = 144'hf4b50c02f35ff6ebfcaaffe0f0a6165915d3;
mem[982] = 144'h029df838f7eb0a341cc3e79a0328ecf8e15a;
mem[983] = 144'hf8ad0451f9f9fe12e88ee19bfcd20b11f7c1;
mem[984] = 144'hfa5b15c506a11d08e448e6261d5a1914f499;
mem[985] = 144'h1084e4fdeddc1bd203a9f17f053fe95bf73b;
mem[986] = 144'he8fd0f0c052913ec1a84194609e31661f313;
mem[987] = 144'h0e16e96af9310fb3f7b4eabd1d89f525012d;
mem[988] = 144'hea280c750dfffa7afffe0d37fbd5ee18e624;
mem[989] = 144'hf92afd07f5d8f7fc066dfd31e2a6f0181b36;
mem[990] = 144'he15405361cdee020f8fde67f01e6f16cfcb1;
mem[991] = 144'h161610d4eea119ccef9c1d81f9cde70dfb0d;
mem[992] = 144'he50717d713f0e045e1671f140734126b1f00;
mem[993] = 144'hea38069d1b9ae298ffe0eedd190ff3a4e9f4;
mem[994] = 144'h025dffa30bc4123df8f61ce7f1081339f32f;
mem[995] = 144'h147419c4fc8614a002e8fee0129a1e550a4e;
mem[996] = 144'hf9e4e0180fa8eae9102414cafb27e1421570;
mem[997] = 144'h1ce8e81316b91569174914481f9708d20b28;
mem[998] = 144'h152c0295ef9402b11dbadfdf1959043709a8;
mem[999] = 144'h07eef0fc0938174be95ee83ff64b0aa2f17a;
mem[1000] = 144'hf169e61be31304141cc70db601b6e769096a;
mem[1001] = 144'hf2811b891021f0271de31e51e7ca1e98f3b4;
mem[1002] = 144'h021402d710c50503f7c1f983e3ec17ce0441;
mem[1003] = 144'h0e8513f1fd1cf470e07a0ee0ef4712c6125c;
mem[1004] = 144'h05f317340ea1efdd1446e32af477e216e599;
mem[1005] = 144'h1d4c1b34168e1984e7d9f7a3eb1a1118fd73;
mem[1006] = 144'hef521ea4021806a012fef926f3f4e1510deb;
mem[1007] = 144'h09d301a0fecbe1c0ee60101d0fd006f617e2;
mem[1008] = 144'hea9215eae923fe110f0bee740eaf1ec6f8e1;
mem[1009] = 144'h1bd0fdf7eb1e1948096119fa1dece075f652;
mem[1010] = 144'h1138e1fff485003dfe5ef630ee8005ff1269;
mem[1011] = 144'hfbb1f5c31c161a54e453fb99e3461064f864;
mem[1012] = 144'hef85130c0e46090deb96ebc00f8f14761956;
mem[1013] = 144'h05c91c42f969e1dce9260f141599ffdd13ea;
mem[1014] = 144'hee32e2be0ac1f22f14fc19c8e107fee30899;
mem[1015] = 144'h0d3ee20df77205a7fe76f652056e1283fe4e;
mem[1016] = 144'hf5a80049fae91c7604de091e16b50de11ed7;
mem[1017] = 144'h141ae0750bb40cee1b6afd021c481f5ff954;
mem[1018] = 144'he075e848f7e51885f22ffd47f6cdeffefc6f;
mem[1019] = 144'h116202ba18ba0ebfe85fec4fe0d7f0181a98;
mem[1020] = 144'h04510a6e1023febf16cdfe4bef75e10cecc3;
mem[1021] = 144'h1c81fd5e1a740da0f553028ef8bce82bf0e3;
mem[1022] = 144'h02a3f4b20f520986ec65f19e0c73077fe5ee;
mem[1023] = 144'h05851003f6201ffe0564f45f051ceb5f0f63;
mem[1024] = 144'h1a7b047d1008134704db198cf0f3e4cf05c9;
mem[1025] = 144'h098ffd66f5e01f271b2bf633f2ba134de2b2;
mem[1026] = 144'h08e514f70feef0b414d2f307e016e638fbf8;
mem[1027] = 144'he5b50a820892e96cfa450cbaf2fc0e41e8b7;
mem[1028] = 144'h17d9f78e16d51269e15ef929f70c0126fc02;
mem[1029] = 144'he80de2850f00e880e625ea29100b1afae4db;
mem[1030] = 144'h094ef58ae2401e7cec2dea5a05a4f28f0df9;
mem[1031] = 144'hef5f08fd20021f27fa530c4218afe4731d7a;
mem[1032] = 144'h0c7c158815ba154c1f8318b7079f09311206;
mem[1033] = 144'h0d34e82e015aee8efa62fb8ef4b2e95fe9df;
mem[1034] = 144'he499e3c6034ce9feee42fea0fd861c271b45;
mem[1035] = 144'hf2e9175117e0086307800197fc0cf6c01395;
mem[1036] = 144'hf23b080dfcbf1c3a12a515fa1afdf4fb0ffe;
mem[1037] = 144'h1eb8f4a91f871c791e3506d81508e27712eb;
mem[1038] = 144'h1acd1d1d009e0362011e0ad81d3ee20c1da4;
mem[1039] = 144'h1119fd81f225f7700164e6e01bdd02be18d0;
mem[1040] = 144'heeb01b8311890e8018dbfdece832fde7058b;
mem[1041] = 144'he778050afdc5e4a2f61102c1e906f29c08f1;
mem[1042] = 144'h1929f0e91fe10ee1f36ff9e2192703cf033c;
mem[1043] = 144'h1bd40e891b7df383ef330b33f168e028e62f;
mem[1044] = 144'hff9de0f81acef7d5e8461a6b08181a34f994;
mem[1045] = 144'hf1690d420906ebebf63712a810faf637048b;
mem[1046] = 144'h0d801334f8bb04c3120915f4f22ff9fb134c;
mem[1047] = 144'h0c58066e0d301c2e11bce5f713f1ef8de682;
mem[1048] = 144'h0e3f09c1f935f155ec08f76710fce462f934;
mem[1049] = 144'he0381fed08e30cf4e4c9fff80e2ffaffea76;
mem[1050] = 144'h1687e6b51a0702d6e366f99bf5ade1411ff3;
mem[1051] = 144'h1f77e8fe1b61199ff2c1fd37e2001cc7e779;
mem[1052] = 144'h1920fde6ee3cec3710991c9aebb1ffc60f0d;
mem[1053] = 144'hec4714f8f53af6c000aaea120f31f9dee3cd;
mem[1054] = 144'he17ee2e017ecef48f7b1ffa10b9918dcef88;
mem[1055] = 144'h120ce087f9e01103009eec9bf39904b80397;
mem[1056] = 144'h109cfee9fc171089f4f004541de3e275f565;
mem[1057] = 144'h09c0fb4e153df4ffe5c105eb1f700ae01e68;
mem[1058] = 144'he3e20b5cf143ea6e1498f358fd06e2c21f1d;
mem[1059] = 144'hf904ee45e40611e9ff4be0711a76ed29f388;
mem[1060] = 144'hfb1c0dc2f137f39f170b02301695e798fc2b;
mem[1061] = 144'he96d10e6175e1cd5e4a9e0e41e73e167e6c7;
mem[1062] = 144'hf564ff1a12000e89fd65feb40f84ffde0b93;
mem[1063] = 144'hec81ec39ec991c9e05b6fff30b9e008a029a;
mem[1064] = 144'h05b507a0fa4cf5981ce0ea8ce5cd1193fd4c;
mem[1065] = 144'hea18f4971c9ff7d61e36e3b915240c3f1697;
mem[1066] = 144'h0698e4681a23f8ca197d1604e288e8ce067e;
mem[1067] = 144'h1df9e4e6f6ccfa9513f71dd002f4fee71da0;
mem[1068] = 144'h013ce5a31b64e42ded8918e8002f1213fd53;
mem[1069] = 144'h0de105e2e3cd0651f49114150841eb13e9f8;
mem[1070] = 144'h163ee3c505eaec69f9a8e9bc1409f2b6032c;
mem[1071] = 144'h1e86045d1b2bf9dff794006b0bdeeeeb0466;
mem[1072] = 144'hffd117bfe5f8f947089b159ff8e80040090a;
mem[1073] = 144'hfd9bef11ea63038bf8faf3e11294e8c60013;
mem[1074] = 144'heb4012cf1ba41af3043410780505107d0c25;
mem[1075] = 144'h05a1038df3a5ff2f1397e50e06c0f0aa14bb;
mem[1076] = 144'h035aedfd0c0b197312fdfce5e7ae1c8ef3d1;
mem[1077] = 144'h0e060ce0f9011fcd02d80e4e188de3180dcb;
mem[1078] = 144'he33ef090f5fc1847e806f43aedd2128af1ba;
mem[1079] = 144'hfc050c071518044aee09e8721fa01768f3af;
mem[1080] = 144'he4310b40f1f8eab80951eb7bfa11f40f0352;
mem[1081] = 144'h0a2ee15fe1a810ebf7d8fc56e402068c1144;
mem[1082] = 144'hf954f70efcf6f8edecc3f5d0f9a6ea8c13e8;
mem[1083] = 144'h1aa8eb9016d9f255ec76054206aaead7e114;
mem[1084] = 144'hf65c0be31f88ecfe156e1c6b0659f5431669;
mem[1085] = 144'hf0ede758e31efe8a0364f164e900141a08c0;
mem[1086] = 144'h1adee77d055f135df420ee741933e330e847;
mem[1087] = 144'hf836f9eeea381873069ee1bafed3f033f6ad;
mem[1088] = 144'h19820d07f8da12ea02a400d6eee70cade9f4;
mem[1089] = 144'h120b19121ccded45ed56ebbbeb3be425119b;
mem[1090] = 144'hf766feee0739f940114c154f19ede547f504;
mem[1091] = 144'he363fa76e0f4f40e19c903c82060ef970955;
mem[1092] = 144'h0253eea0f78a1b4cff7e1d87e401f68f1f47;
mem[1093] = 144'h12e0e518fcb11513eb3011851ee2f5d60108;
mem[1094] = 144'he194f5641bd601a4f605ec8af6bd0b61eb52;
mem[1095] = 144'hed69f812f23af4d8f2dd087deadfe808f01e;
mem[1096] = 144'h15ec112dec83f1570f7e0986e6b50bee1623;
mem[1097] = 144'h181eec2d1015f2af06c9f293ed32055417e8;
mem[1098] = 144'he987e669e7291e5cf25b0bc20606f82ef350;
mem[1099] = 144'hedd01393f2a20b000372f6161c40000bfc6b;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule