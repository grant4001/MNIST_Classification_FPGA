/*
Copyright 2019, Grant Yu

This program is free software: you can redistribute it and/or modify
it under the terms of the GNU General Public License as published by
the Free Software Foundation, either version 3 of the License, or
(at your option) any later version.

This program is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of
MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
GNU General Public License for more details.

You should have received a copy of the GNU General Public License
along with this program.  If not, see <https://www.gnu.org/licenses/>.
*/

`timescale 1ns/1ns

module wt_fc1_mem6 #(parameter ADDR_WIDTH = 10, DATA_WIDTH = 144, DEPTH = 1024) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h06e2f21100060525f2af0229f2a3031d0c30;
mem[1] = 144'h0704fd7ef9adfecb0aa905350d700b1a0f35;
mem[2] = 144'hf9caf01d0148098a07b4f95707d5063afec8;
mem[3] = 144'h0da6f3cef85f0dfb06e5fa5c0f9e03c302f7;
mem[4] = 144'hf7bcf841f6d8f98efe97f03cfca30691087c;
mem[5] = 144'h096bf56502f1fba1f9a7f507f1230a680829;
mem[6] = 144'hffc1f6010caef5d308a20304f915f73d0f93;
mem[7] = 144'hfeb5f93a03b8f26a0b9ff8f305eff7c60829;
mem[8] = 144'h05cffebafb720baffce70e9d0e9ff6fbfeb4;
mem[9] = 144'h02b40107f967f6b1017d035cff5af04b05d1;
mem[10] = 144'hf0baf15df45b0b5efc530d0ff8490f0df2cc;
mem[11] = 144'h0c10f2d50c000aa9f562003e09d8fd8606c9;
mem[12] = 144'h08f707a300e60242f127fc65f6cbf40a04ea;
mem[13] = 144'hf9a50b710e9a0d1603ef0ce0fde10ea20a28;
mem[14] = 144'hfcfbf311056c016dff71f802f0aef4b2f31b;
mem[15] = 144'h0e1f0448008df7e1f40c0abff7960ccef784;
mem[16] = 144'h0fd5fae0ff73f1e80f4dfe0df69ff0bf0540;
mem[17] = 144'h090a052af948040704edfde4fbf007b9f96c;
mem[18] = 144'hfaa00818f53c0046f88ffdf30ba502c50c1c;
mem[19] = 144'hfd5efc46f7e6013800abf651fc47f925f1c6;
mem[20] = 144'hf395098ef930f7ea09a2fb9bf5bd0caafe2b;
mem[21] = 144'hf692f11cfbca0df7fbc60ec301d4f1d2fbaf;
mem[22] = 144'h0aa10033f35af7a0fe80fa15ff2afe8c035e;
mem[23] = 144'hf73e075df7830fa3f10cfe54fba4f13e0509;
mem[24] = 144'hf55806550abefe9ff16ef945f25000d8ffff;
mem[25] = 144'h0b13f005f57d042e0014044a043a04150d35;
mem[26] = 144'h08df077ef248ffc1f788f0d40f7bfbd1f273;
mem[27] = 144'h055dfdcb0d9effff084bf21f0e58f2d50ae8;
mem[28] = 144'hfbccf0d4f9dd0359f309f70703a4f78d0b5d;
mem[29] = 144'h03a80b0cf06c0fabfe09fadef77ff3c7081c;
mem[30] = 144'hf92d0bb60e3bfbdbfd13f7420d69f2d50586;
mem[31] = 144'hf8500719fada0c09f89f083c0a630d2df999;
mem[32] = 144'he3a2ead7f5e0e68bffbdf0a5f64ff378e09c;
mem[33] = 144'h0d9ff998faf2fec80b30f0920f8c04f20b4c;
mem[34] = 144'h0c9503e908fdf160f7130506efe30a3103dd;
mem[35] = 144'h039b036d061ef4e6fa2cedcef39ee086e9d2;
mem[36] = 144'hff0bf80c040def19f23004e40946ee9ff0d8;
mem[37] = 144'h02670a87ff2afe16fdd7fe6a0c99fa15f3a1;
mem[38] = 144'h074ef64200f907b900330c1ffe110d9c0d37;
mem[39] = 144'h0d7a0681030fef49067c0ba5042cfa86f055;
mem[40] = 144'hf7d6f95a0c99ffb10a8b0bd3f3dd0286f6df;
mem[41] = 144'hf79bfcd0f00b06a90a1bfc4e08ecf5b3fa2a;
mem[42] = 144'hf1ea02b90f5b0916ff10fe15fb090f710244;
mem[43] = 144'h0bfd0bfafe3606770848f2170815027b05dd;
mem[44] = 144'hf6ebf8ddf720f6e3f301030af9eafcd2f5b2;
mem[45] = 144'h0daa09a5fd570aaafadcf487092bfff5fc24;
mem[46] = 144'hee67ece7f4a9f447e479f612ea51e963f02b;
mem[47] = 144'h0120f5effbc9ea28ec94fcf8f1c9f9a9eee3;
mem[48] = 144'hf48eedeaf304ec02f765f159fdfee0ebef83;
mem[49] = 144'hf165028bff0a08920aeffe0f00cdf1e6f33d;
mem[50] = 144'hfe75fa0eff4d0a2ef3e8f7300a890dc20124;
mem[51] = 144'hfb84ec7de808ee5afba902ef0423030ff7d8;
mem[52] = 144'h0b9503290944f400f97bfae40a2ffae20cbc;
mem[53] = 144'h04960dcbf71cfa7e0c3af177053cfeb8fda2;
mem[54] = 144'hffecff5ff759ef3f0da50e760e5b09f50bb4;
mem[55] = 144'h03010e27f79307ce049e085a01f80417f2e2;
mem[56] = 144'h00b0030ef46a0dc208adf2e1ee8b04cc0ae9;
mem[57] = 144'hfcd3f1b1f7e2f36df5e1f566049a093a0bb1;
mem[58] = 144'hf363fba204b80d8a0874e320f4d5f3280742;
mem[59] = 144'h016e0aef0234f315f2c0fcec0b90f8cef098;
mem[60] = 144'hf01bef6bfbeef426054605440f57edd70746;
mem[61] = 144'h0b89f21ef680f3b2f8de07890b3cf51efa02;
mem[62] = 144'h0b71efb6013aeb46fbc3fd780248058504dd;
mem[63] = 144'hf03ef5c3016ef3f0efe4f49ef1ac081ffe5b;
mem[64] = 144'heb0df819029bfe230721f730071dff65f789;
mem[65] = 144'h08d9f437f282054c0717fd7701c609d0ef07;
mem[66] = 144'hef1b031b08b7f39c02160b6c094e09c9f1ec;
mem[67] = 144'h04f0eeefe91efeda02d1087dff04f267e24a;
mem[68] = 144'h06060b490606f700084ef5cdfe72061c0135;
mem[69] = 144'hf20b00e2f42100b304540a720d400862023c;
mem[70] = 144'h0eedfcfe05c8f02ff4390cf90299fc61f148;
mem[71] = 144'h0997f0c60baaf21c0944eeafefd906ad0804;
mem[72] = 144'hfc08fb4c044bee0cfe4d07de0ab007d3ffba;
mem[73] = 144'h06910383036df0c1f94ef4b1f5c9f9450af9;
mem[74] = 144'h0017ebbb1752079df58ef57cf849f2ca0fad;
mem[75] = 144'h0e2207d2f94703ee05f9f1f8fa49fe44f6fb;
mem[76] = 144'h034e03a206c707b5fc2afc72fe5be98cef2f;
mem[77] = 144'hf0a905d8f9b8ff1cf1caf266f299fe4a0256;
mem[78] = 144'hfa84f20ef534f564fb170420eddedc14ee29;
mem[79] = 144'hfcf706dd07b2f9d5f575ee5a0325f0bff7d1;
mem[80] = 144'h060cf545ec3aea3bf082f3e2ef3ffacef682;
mem[81] = 144'hfeb0f5fff39801d7f52df04bf590fe690afc;
mem[82] = 144'h06f2f20f0e3df8e00380011f0107fa11f04d;
mem[83] = 144'hef5e0450fccdebf305fef85609fcfba2f216;
mem[84] = 144'hf238032701500d6ffb910e56f61500c3fc6e;
mem[85] = 144'h06b6fad809d5f1150872f0990bed0c09f97b;
mem[86] = 144'hf1adeff803bd09d305cdfb37ffa1067ff8ba;
mem[87] = 144'hf48509f3059f0df0f713f0daf2def1ddfca3;
mem[88] = 144'hf32aee530e73f9fbf659f1bd0af90ad50740;
mem[89] = 144'h0971061ff2def5ad049a09cefe8402e8f2e3;
mem[90] = 144'hfbeef6dbf70207cf0227f0ebf130f4fb00ef;
mem[91] = 144'hfbbaf06c0358f03bfdc9051a0c6ff990f059;
mem[92] = 144'h07530628f423f862f61d00fa0ad30d69fe05;
mem[93] = 144'hf88bfa8309c10b920963023efec10f15fa00;
mem[94] = 144'h0c3dfac8f2bbf21d034af38df5f9fd3f0785;
mem[95] = 144'hf349fc6f04230c2f06f901a00940f45205c2;
mem[96] = 144'h0a6ef6b3051cfe01074d03e0f49df2240440;
mem[97] = 144'hf7d8f696f706f451f22802c9f63e04c60b06;
mem[98] = 144'hfbcd09c40925f8fc0d6a0d28fcf90459f1f5;
mem[99] = 144'h0e51f18c01b7f1dff40ef08f0d6b04ed00dd;
mem[100] = 144'hf4a4f1b20e680dd70ec3f7210d390959f3d7;
mem[101] = 144'h0de70bb1fd8afbfc03d60bd3018fffe30eb7;
mem[102] = 144'hf33df5b3fe48f402fb23f3d3f6fbf057f12a;
mem[103] = 144'h0205020efe0c089f0921004c0a42f40efacb;
mem[104] = 144'h0a4f0d1e0e3501c00d57ef7bf0260aba03d2;
mem[105] = 144'hf83b0a63073af178fd230835f9a6f0e2ff39;
mem[106] = 144'h018a06b3edf40230078af3400a12fb43f6e7;
mem[107] = 144'hffcc0bbd017303bcf202f154054b03eef16f;
mem[108] = 144'hf178f7baf9020d7405640f680963074d0dec;
mem[109] = 144'h0718ff10fef30027fff90351f8640f1305e4;
mem[110] = 144'h078af24900b6f402f4520cb7f61ffb870a69;
mem[111] = 144'hf01703b60800fe86f12801180dfd079108fd;
mem[112] = 144'hf1a6e7b502b7ef890b6bff07fc14f526fd59;
mem[113] = 144'hf08c053cf3170322ffb7f953fef30c46fa00;
mem[114] = 144'hef51fa0ffebf095a0dabfeac02310b5dfc9b;
mem[115] = 144'hf06a06cbf0e20701ef7008090cadf976fd41;
mem[116] = 144'hf810fec0047cfde7f7ebef5ff3f0efa8f689;
mem[117] = 144'h062601a100590594ef54091c0423fc4d0a5e;
mem[118] = 144'h077b07420715f89af0daf71a0469098ff314;
mem[119] = 144'h0685f907f968f0b305a5ff35f3a409cd067d;
mem[120] = 144'hfe3606b0f11d0608f1f5f8bbeeb7fecef2cc;
mem[121] = 144'h03e4fbf1f673f4c0fef30245f09b0218ef98;
mem[122] = 144'h087ee15116a7feb4f2a1eee706dbe9ef0582;
mem[123] = 144'hf517f73deeedff51f0cc047d09cceeb3087f;
mem[124] = 144'hf2050cc60280f533029b036cf7bb081a0a0d;
mem[125] = 144'hf351f68006b606b10cf0f4cd0d11fc1a040d;
mem[126] = 144'h0c8fed0bf0ef00f6f937f8b8072008a8ea57;
mem[127] = 144'h0af1ee6beb5b026a00fb0794010300ecefaa;
mem[128] = 144'h0094f6f902b5091b03b7f37cfa62fdb2f1cd;
mem[129] = 144'h092ff80af2ef0d96f2f80a66f6fcf37df320;
mem[130] = 144'h0465f33b0bf0f52509a8fbf0fab405e7f605;
mem[131] = 144'hf563086300a8f204fcfcfc2a0cd7f589fb5a;
mem[132] = 144'hf2b608bff66302c50897f85e056a0f3f00fe;
mem[133] = 144'hf691fef105ea01a6f1f5fc510af400430e23;
mem[134] = 144'hf2edfa20fab3f672f965ff64fade0da307e6;
mem[135] = 144'hf3ec0a6b085c0be90998f772f39a0cb20989;
mem[136] = 144'hfc3a0bb8f23df9fb0484f774fa61f58af39b;
mem[137] = 144'h032bf137051701ef0539f9d6fa140f59ff02;
mem[138] = 144'h07130169f0eaf1cb015800caf3b5f097012f;
mem[139] = 144'h076ff5dff073fa76fca1f78005220be5f1c9;
mem[140] = 144'h03daf7e5093ef82ff0aaf3980acff99cf16d;
mem[141] = 144'hf9baf4ab085b0e6a073b027e0b6d065502fa;
mem[142] = 144'h01e70f27f5ff080dff2803b2fb61fc1afd97;
mem[143] = 144'h027f0b77fda2048dfbf10478044df7970e9c;
mem[144] = 144'h009509a209cefc5a06a3fd8bf2a804d5f683;
mem[145] = 144'h0bdef880f5dc0f38fd8d0d2f0d49030a0400;
mem[146] = 144'hfd47f2eef88a070b0352062b082d0f8af252;
mem[147] = 144'h000308c5f5cb0718f4faf3fdf0c00dd500ba;
mem[148] = 144'h07b8ff65f44906df048f09b1feb3068afd66;
mem[149] = 144'hf4e40b8108bdf41bf5ba0444058e0d3d0dc5;
mem[150] = 144'h040afa93f484f57407bb0d1505c4f08afc1b;
mem[151] = 144'h0ee2f843f9390b57f229fb06ffea0b9cfc3f;
mem[152] = 144'hf65c0ad1feaef9edfc61fe12094300bbf955;
mem[153] = 144'h0bcbffbff9af053f001103420e1df110feef;
mem[154] = 144'hf87207bdf4f10cb004d1f92403a30008f153;
mem[155] = 144'hfcf4040101b6fdb1ef90030e041801e60389;
mem[156] = 144'hfef50c190bf0f7c70f93fe0efe3cf4ab06e6;
mem[157] = 144'h07e1fd50f40cfc65060d0fa0f4b0f92bf661;
mem[158] = 144'h0863061ef98607d9005dff0b04caef770849;
mem[159] = 144'hf6a70bd2fc29ffdbfa0206f10e73fc80f13d;
mem[160] = 144'h05aafb390d76f78efec50cdc09b8f6b6f526;
mem[161] = 144'h08cfff5d05db0722f9f4f88ef8dff07ffcca;
mem[162] = 144'h02edf34f0e1809c40c6c0832f311ffd1fa51;
mem[163] = 144'h08c20c0e0103fcb4f5760443f2b0f046f213;
mem[164] = 144'h005bf1b5f6120f62f45409600aef0ed40c5a;
mem[165] = 144'h0d04f567094df60b006efadcf522f1e3f07c;
mem[166] = 144'hff64058003f6f5db091df8e20ccdfe3a065f;
mem[167] = 144'hf22ef2e30e07fe75043e051ffd51f888fc0f;
mem[168] = 144'h026700920566f5dbf0b4f8a201000c8dfa9e;
mem[169] = 144'h076bff32f7f6f7440750fe72f7b1f344f06c;
mem[170] = 144'hf912011d0bd5ee9f0872f4caff41fba100df;
mem[171] = 144'h002d0987f5f1fd0cf2010331fd6b0aad07e0;
mem[172] = 144'hfe07ff1bf118f4fff61f09defcee0188f849;
mem[173] = 144'h0e68086b037ff585f46bf3b10d2cf633ff36;
mem[174] = 144'hf1b800e10db5f58dfd1bfbc2f17efe3af8b5;
mem[175] = 144'h06c50e800753f34f027101ba0208f4ac08e3;
mem[176] = 144'hf986050f03d8f264082d0216fcc7f2830d75;
mem[177] = 144'h0ab1f6f4014cf5f6fc1cf96d0e76f2e10da1;
mem[178] = 144'h03aa03a80f8e07b8009a0d12fe6cf8b0f72d;
mem[179] = 144'hfb540bf0fad4f392f3def0fffb6e021bf885;
mem[180] = 144'hf53a0523f30c0e00f2ddf408f0bdfaecf496;
mem[181] = 144'hf878093e0d640dccf2b5f6f0f46bf4ddfe4a;
mem[182] = 144'hff6f030df8a40e6906b10445fa3d09cdf2aa;
mem[183] = 144'hf637027fff4af0f70c14f3f905f80379f762;
mem[184] = 144'hfeea04b6f351f4250149f1f20e9501740708;
mem[185] = 144'hfddc038ef6fe0ebe0b22034202560452f3a4;
mem[186] = 144'hf640f0af08860eb7f971034f0ca9f6a4f42f;
mem[187] = 144'hff410672fd33f2990f8bfc0a041905c40707;
mem[188] = 144'h0bfefb72065ef1a6f68af1a5fcd9fda60dfd;
mem[189] = 144'hf7fe0d64f70eff72f962f18cf1a7f829f789;
mem[190] = 144'h07b80ce3f369069cfa010528f16906260f58;
mem[191] = 144'h0daa08af0d62fa840f01f672f1daf513f8cc;
mem[192] = 144'h02490d83f01eed7aef54071004eafed0fe54;
mem[193] = 144'hfa83fb43004c0a820f9af2dc09e00ced0b54;
mem[194] = 144'hfd8ff58d0cc308b1feaff1f4081405f0fa8f;
mem[195] = 144'hf88eef1ffe9fee9c0759f0dff2e20f1efdbe;
mem[196] = 144'h0227fc99021fee130d82f32cfe3a02c3fe18;
mem[197] = 144'hf4cd0bd5050e066d01320ad1fa5e07ef04d2;
mem[198] = 144'hfd53fc97f0180198f2dc02bcf984f20904e3;
mem[199] = 144'hf69906d604dcf393f82fff1c067709a3f9b3;
mem[200] = 144'hff91f333f09cf3d3f81d0a42f317f9be0791;
mem[201] = 144'h0b2c0c2d00b4f4f90c3903db0d26f9d70f0c;
mem[202] = 144'hfe550405ef93f68d06a6fd7c07ccf04ff1fe;
mem[203] = 144'h07c00a8009c1f8e1f77f0d97f2e5f611f198;
mem[204] = 144'hfa7af1fe06ae0ae1f49b03b60c16f49403ab;
mem[205] = 144'hf849f92e010302450405f084053704f9fe77;
mem[206] = 144'hf8dbf3e0086801b9f601f862f12af0f4f235;
mem[207] = 144'hfc58f491fecc059908d60c94f085046ffd4c;
mem[208] = 144'hee17f240e69108cdf3950eaafff3ff8cf6bd;
mem[209] = 144'hf3c4024c0cb2f2350a8005abf91900670329;
mem[210] = 144'hf02cfb40ee81043ff6ea08da01ff0d900003;
mem[211] = 144'hf208fbbcf2c605a00546fadcfa23ee05f243;
mem[212] = 144'hf427ee20049e08aaf132f06efac4fc1b03a5;
mem[213] = 144'hfbdf06ba050f06f601cdf13f076a036909c9;
mem[214] = 144'h023108c00e3b0721fbfefd5ff23cf8d4faa4;
mem[215] = 144'hf8cff5f1f7f60c65f585f06d0cd405d3fee6;
mem[216] = 144'hfe7e0316f2b8f7180b0e0b1208a00026fcae;
mem[217] = 144'hfcf105f5fe2502d2ef3f0621f5fef54e02a0;
mem[218] = 144'hfa7af474e1560fa00b11ec27e985e3d7fa58;
mem[219] = 144'h0078f31708b0f227f906ed0cf2e7ee790b2e;
mem[220] = 144'h01eafa4af152f7f60a200bddfdd2f675f204;
mem[221] = 144'h08d6f963006ef90b0cf4f9ec010a07b00cc1;
mem[222] = 144'hee42eae5f3d7f775f52afdf30065eaacf79b;
mem[223] = 144'hfba4f03804acfd690caa0e13094408fcf824;
mem[224] = 144'hfc2beef9d6c0e17fefa202b0ea89eee3f80b;
mem[225] = 144'hfb49071f03d606c20da906b3ef4003690bbb;
mem[226] = 144'h06b3098b0267086107b4f539ef5df63a0e69;
mem[227] = 144'h0a70ffcb00b4ecd3fdf3057205a4fa4ff4ee;
mem[228] = 144'hf22f019cf828f4ebf89f084bf038094e0334;
mem[229] = 144'h0b7607e4f37f0042f9440bc6ef0a0447f28c;
mem[230] = 144'h07ed05daf3920ad90d0b0a81f678f668fd5b;
mem[231] = 144'hfff0fbeafbb4ff1d00a8eeeafc30f5c10cf2;
mem[232] = 144'hf9ea071b0993f6ef0642f1ab0559fd660606;
mem[233] = 144'h09e70ecbf890f165fe88f0dbf472f8fbf203;
mem[234] = 144'hfbe10c050eb1177bf677fa97e3fff248e9ae;
mem[235] = 144'hfbebefc6fd3af116f77c04fcfca8faf4ef9c;
mem[236] = 144'hfcb2ff7ef4c5f29cf1dfee540a0808aaf722;
mem[237] = 144'h09610686fa770ecafd420364ff050ab30221;
mem[238] = 144'hee28f0730502f0dbeeaafe9f039eeea4ee65;
mem[239] = 144'h0237f778f90908b7f2d5f7e30a69fd4df320;
mem[240] = 144'h060b0df00cfb0e2ef4e3ffc4048c0c02f1ce;
mem[241] = 144'hf7e0ff5706a7f172f7fd03cffa8bf717f626;
mem[242] = 144'h0734f9fcfd2dfb4602ff0a98f020fcadf68d;
mem[243] = 144'hf836f1380c13fa35f35df47c0b78fc21ff2a;
mem[244] = 144'h02affdabf4f4f1fdf4a502860d42f1bc0922;
mem[245] = 144'hf55802440b46052904bb04e5f7280503f9a3;
mem[246] = 144'hf3330e59f6dbff06fd55f37a0ee60be108df;
mem[247] = 144'hfbd1014cfffa0cfa098cf69c009cfea5fa41;
mem[248] = 144'hf339ff0df51205dff08d088009a5f6740973;
mem[249] = 144'hf39a009cf696fbae008cfe1805fafa6208b2;
mem[250] = 144'hfbefedd00a4407fff306f48ef3b102f8f1a3;
mem[251] = 144'h07fb0645f8400b4ef36900a6f694fa75fec1;
mem[252] = 144'h01b7fad30138f26a014ff6060148080afe84;
mem[253] = 144'hf2c30295fc8303affcd10e78f501f26ff230;
mem[254] = 144'hf8aa0825010af3b601a405c00ed8076708ae;
mem[255] = 144'h04c8f8a408400c79f0a4f1a20d9d0d2d0a4d;
mem[256] = 144'hfe1af83ffe21f9e70dbf0094fa11f767f600;
mem[257] = 144'heffe02c7fd41043ff16bfbd7fbfd033df7d8;
mem[258] = 144'hfc4df809f1370d1af027f41ffe1ef401fbdc;
mem[259] = 144'hfa51f5970735efd60342f272fa0e0d27fa64;
mem[260] = 144'hf8b60d5a0b980b460823fa950e80fe78054c;
mem[261] = 144'h06170ae3fd01fb81fc4cf57ff075fa7af754;
mem[262] = 144'hfeec0bd3f2bbf04bf364fed3048007eaf8f1;
mem[263] = 144'h0dd50df7f344f05406390409062f0c990cb2;
mem[264] = 144'hf9800b82f980ffe7f3e20969088f0f640db1;
mem[265] = 144'hfa580ebffc1affa5f6a20e58f08506cc026c;
mem[266] = 144'hf9acf56f08d804c8fd8ffb17051af3ae05c2;
mem[267] = 144'hf5ce078ffcdeee53fc63f67606abef1e0ac7;
mem[268] = 144'h04c6047efb2d0e9cfffb0aaf08dbfe4c0740;
mem[269] = 144'h0280f2b1fb6e06940a97f7b1fe84f566fbc3;
mem[270] = 144'h00baf97108ff0418faf7f64bf657f325ff6f;
mem[271] = 144'hf880eea6017cfd51f7d106ef0ce0ffd202ef;
mem[272] = 144'hf50a053d095f0eaa0b210365f882f708f90d;
mem[273] = 144'hf961fa30f7e3f1e50a92042cf2fbf286f011;
mem[274] = 144'hf1a30a2d0d9301b304e6ffbef716f7fb0fab;
mem[275] = 144'hf195fe8df3330286f621f06a0cedffb5f4b8;
mem[276] = 144'hff7cfc55f3ab0cb8081c0839f78cf6a20147;
mem[277] = 144'h086ef0dc0cf706990b07039105a8f110f740;
mem[278] = 144'hf37c03900f16fa55f8bbfa79fd1bf90dfc43;
mem[279] = 144'hfa9f0da30081f9d5f5dd02380c690371fb93;
mem[280] = 144'hf215f4eefcaa0995028d0e3bfe120fb5040b;
mem[281] = 144'h04dc0e5b0909f048f8f4fcec0608f236fa36;
mem[282] = 144'h0d4bfc0bf63c0d73fc80f9b307e4fd0200ec;
mem[283] = 144'hf7cbf882f13503d20f9ff61ef6def4ff0388;
mem[284] = 144'h02db01730037f2400cb6048af4c902760af7;
mem[285] = 144'hfc2efffbf5b600b7f396025df86df09b0e19;
mem[286] = 144'h0809faf4f730081403f7fea1faacf025f9db;
mem[287] = 144'hf91e0c3efb17fc76f4630e0dfc1ef7c6fa78;
mem[288] = 144'hf657ee88f850f282f24e084cf6c3e92a01e8;
mem[289] = 144'hf6e3f94c0d370bde054e00590d8503fbf191;
mem[290] = 144'h0d9af510064f09e20ced0a13fb27fc09fdc2;
mem[291] = 144'hf3fff289f8b1f056f34cfec80238fbb20070;
mem[292] = 144'hf277f3c50d20f675f1c604c5f9550361f11d;
mem[293] = 144'hf67ff5b7ff8903e4ef240ebe0962096c0030;
mem[294] = 144'hf42d0e56f45ef5ea045cf5d4f715fe5e0b9e;
mem[295] = 144'h046207ccfbed0af20a33007e0efbfa34ff61;
mem[296] = 144'hf3b70487032bfbd900b7f449072406d1ef33;
mem[297] = 144'h08eefa31ff8feff7f3ddfed20c1cff7af428;
mem[298] = 144'hefc90d070cc9072e11b7f9a3ed57f52c0d68;
mem[299] = 144'h06ad0103efbcff6e0150fe54f0320603fa84;
mem[300] = 144'h0b0ff118ecf50c80053ae99901fb0b3ff08d;
mem[301] = 144'h095506c8fd710411fb88ffc70c93f32a0f28;
mem[302] = 144'hf282fbccece8e225e969fd8bff83fee0f600;
mem[303] = 144'hef8305cff21bf35f0708feca099df379fe76;
mem[304] = 144'hfdf7fbbbef24e34501d602e8fd22f8bbe489;
mem[305] = 144'hf536f3c608adf40e028d048bf4acf4ba01dc;
mem[306] = 144'h0b1e03f6f19b0e11ff58022cfd3bf90e0ddd;
mem[307] = 144'hfeba0626efaeec4f073b03f8fc02f52df491;
mem[308] = 144'hf09df27ef31a05660aa3f734040705d6fb9c;
mem[309] = 144'hf7ef0be3f3dff0b8067afa3107d0eeaffe4d;
mem[310] = 144'hfaa2fe3705c00b6a0a5a09b303b8076d0c42;
mem[311] = 144'h08abf4aa0698f0a4055defc9fcaf0d28f53d;
mem[312] = 144'hf72ff2d4fb63f9f507730ca60c9f06bef1b1;
mem[313] = 144'h05760751021bf230f44ffcc8f5bcf2330517;
mem[314] = 144'hf1f2e916eec30d1c01a0f83bfcd00618ebe0;
mem[315] = 144'hfa1ef369fb4b027509080536fa19f708fca9;
mem[316] = 144'hf0c3f5a9f7daf1a20c09ef890f9af6fc0076;
mem[317] = 144'h0afefe7b0ae9f7a0fca6ff9e04f70c1cfc7e;
mem[318] = 144'h0bc2fd19fb4ff197f349edf4040f0285f39c;
mem[319] = 144'hfa5bf8890c4c0af6f79fef4c01600aa50966;
mem[320] = 144'heaf7ec09f251f384e38c0674f835f100e6a1;
mem[321] = 144'hf93a09f507d7f0d9f5fc0bb2f275022df82e;
mem[322] = 144'h08f3003b05bb09040186f7b9f0350bf3fe30;
mem[323] = 144'hf48fe453e9dee15de4d0fb2a0788eeebf4b8;
mem[324] = 144'hf4e4fc5209edf91bf9f4014ff618eec4fb5e;
mem[325] = 144'h0be9018c0a0807f5080dfc7000160992f687;
mem[326] = 144'hf2a70205f336fb84fad209fc0b39f8fd0859;
mem[327] = 144'hf0d6fee00bc20df0f0ed0192f8f6f74805f0;
mem[328] = 144'hf26dfff5009df542f5280b00f31605c0068a;
mem[329] = 144'hf96902cbfc1cf96dfb97fc8af553fe10f7ee;
mem[330] = 144'he7a7fc110389feb906ecf6bdeba3f2790992;
mem[331] = 144'hfe1c01c5077c0c1bf7c9f02ef83f02b90900;
mem[332] = 144'h09b4f10cf5aff143e42de7cc0495f996fcc0;
mem[333] = 144'h059d06cff21908a100eef500f4c4f3c9f313;
mem[334] = 144'hf237f822e40cfb15fc09ec330861f319ea49;
mem[335] = 144'h03ffffe1ffb202abf303047df3a4fb8901f2;
mem[336] = 144'h0695e95a05a0fa10f21bfd27fd3800f7fc36;
mem[337] = 144'hffddf8c2f168f879006bfa5bfeda0ea207bb;
mem[338] = 144'hfd3e010ef82ffb57064bfb46faa0fdcb0e44;
mem[339] = 144'h003eef2feb10f60ffd18f47c0c5408a7fce1;
mem[340] = 144'hf3f6f94a030b0345faddfdcb0c33faba03a8;
mem[341] = 144'hf4c4fe4006a2f75df10cfec7f6a3f9780cd0;
mem[342] = 144'h0ccdfb4c0628f9f00d8307650c58f86bf900;
mem[343] = 144'hf14bf5ddfd57ff260b9802bdf4a8f6030852;
mem[344] = 144'h0b1a0c67f4e309eefe440592092902ddf7a1;
mem[345] = 144'hff9e06a20585f5d9f64c0c66065b06320663;
mem[346] = 144'h051ce6fd003bf5d6de4d098cf5e701f103b6;
mem[347] = 144'hfbe2fb6ff87009c2f1390d36f51bf3d1f1c4;
mem[348] = 144'h0e47017802f0001c078def7a0663fefa0904;
mem[349] = 144'h08b10d040facf4090fd8f6830025042604a5;
mem[350] = 144'hfa94f4bcfdd6ed650632fe48f03309f8f8a8;
mem[351] = 144'hf291073aeceaf93307eaf86a0d33fcf40aa4;
mem[352] = 144'hf13f0149faee0467f55b04b0e7aafccbeda1;
mem[353] = 144'hf3d90c9c0c9004bcf1c401d5ffaa04e803bc;
mem[354] = 144'h0c4df9f90e6a02d5f1940107fbea00a000bf;
mem[355] = 144'h0800ef89f45102f9fbfe00f1f692f7fef487;
mem[356] = 144'h0908f15ef430edfb03b5f56ef3e70a92fe8f;
mem[357] = 144'hfb05021106bbf1a70d8df1a50b73f5980da2;
mem[358] = 144'h052209a50d010176f4e5094a033f0b3af084;
mem[359] = 144'hf1c6054e0e620c0400b50137fbb2fe51f191;
mem[360] = 144'hf394f13dfa3ef0600151fe6af906f31d0a96;
mem[361] = 144'h04700105fe05fa4c0b45f9c2fe34072c0e3c;
mem[362] = 144'hf55deb030fc8f5a9ec70f46dffb50d3f0443;
mem[363] = 144'h00c70deafcf5f34eff9ffd8ff6e5fc02f40b;
mem[364] = 144'h01cbff32f9c7f605ed0ef4620198ee8e038d;
mem[365] = 144'hfc95036000e30480029bff08008104a4fc4b;
mem[366] = 144'h0045f8adeb54f9c1f6a003e9edc4eecbffb1;
mem[367] = 144'hf194efbf00860a0f0174fa20092cf88cfee4;
mem[368] = 144'hf800ffa703b4f62d0479f5a00948050005fa;
mem[369] = 144'hf626f37e04c4f67cfda4f0def19afa86f595;
mem[370] = 144'h0b4ef48bf49a00b2f5d30e02f999fffcf42c;
mem[371] = 144'hfc2ff7fbf912f8720793f156ff510a1a0262;
mem[372] = 144'h062af6bff43b0a9af37902b90695fd5ff6b2;
mem[373] = 144'h0546ffbcf7210b9bfd4b01a30a9afb46f650;
mem[374] = 144'h02a5fd1b0773f66f09f50dc9052301d7f51e;
mem[375] = 144'hfbdf0b6fffa201f200b00b0e06cb063a0d6b;
mem[376] = 144'h0dbe0cd4fc3cf9bbfa91efe3f8840cf609cb;
mem[377] = 144'hfe4607ae0929f91cf91201c90fcaf826f6af;
mem[378] = 144'h0e680502f4260c95ef7ff3c70363f1f5f95a;
mem[379] = 144'h0ddbfd4ef8a4fd93f173042fff8e0c410be4;
mem[380] = 144'hf41ffe7e0196f9400cbc0fd00e0d0f59eff6;
mem[381] = 144'h07e7f230001b0fdf0ff1fcea0a1af4c505f4;
mem[382] = 144'hf4f6f75afc0cf383f5750f7ff28af9220f95;
mem[383] = 144'hf29b0ba1f34a03a1070cfe58f0630434f124;
mem[384] = 144'h0d99f5abf90008b50b220bccf899fde90a7b;
mem[385] = 144'hff88035c0e2f0f06f60df6f4fba8fe5af8f0;
mem[386] = 144'h049ff3d102f903630c14f9100d42098afab1;
mem[387] = 144'h08cbf146022004b4f6d6f30e0391ff5f061d;
mem[388] = 144'hfacd02e30676090701880b65f31bf73bfed6;
mem[389] = 144'hfbc802e3f3c5020100c2fe350d94020ef485;
mem[390] = 144'hf4d4f84bf6f8f2f306130991fe2afbd8f7c5;
mem[391] = 144'h03f5ffa7f6130654f9b9095503aef25408c6;
mem[392] = 144'h0a97f227ff91f4250be0f1510a25f83af5db;
mem[393] = 144'h03def11ef66208fdf371f24bfc8201500854;
mem[394] = 144'hee82099c0154f8e7fa4a081408b1f8b3edeb;
mem[395] = 144'h0eaff6950ea7fa3bf03efad104fdfa8c0491;
mem[396] = 144'h08d1f86bff590a520b18ff41f5c0fc6f0994;
mem[397] = 144'h011cfe2df74604fc0286fdb7f96509ddfb7d;
mem[398] = 144'h0d85f82bfc64f908f26bf83a0155f525fa9e;
mem[399] = 144'h039a0d8b0ac80906fa16087cfd330639f848;
mem[400] = 144'h00edd81ee901e84e09d2f7cc01d6e9baf68a;
mem[401] = 144'hfc8ff8020044f011fa2d08e40122eeb6f33c;
mem[402] = 144'hffc409bcfde9f4ed0806043cfe3f081b05d4;
mem[403] = 144'h04e3fa4be92af8c2f895f53bfa93fa47febd;
mem[404] = 144'h0220f6f6eebef7890bb406b6f7c9f466ef82;
mem[405] = 144'h03deeff0067801c7fdb9f51b0b0dfb74fc40;
mem[406] = 144'h02b3f76af641f85903dc06e9f486f25ffe1f;
mem[407] = 144'h0a41fdb4fe2c0bc805e90b5cf857ee92ffd6;
mem[408] = 144'hfe54fccd07730142f557f610f6790bfe0938;
mem[409] = 144'hf9150367098d0dd4082f0dc50ad70eea001c;
mem[410] = 144'heb210127f0da011e0a93f2400056fc16f8c4;
mem[411] = 144'h04560755f6f70e1ff79aeee9f75a0d78f586;
mem[412] = 144'h0ef8f357ea37031ff067fa86008dfd13eec4;
mem[413] = 144'h0a06fcef06fffd730dbf083ff06c0616f4a2;
mem[414] = 144'hf464f5bde493f61df9a0f1b3f3b8eb50ee42;
mem[415] = 144'h023af1c6001e04a2ee8e05d308c6f2c8ec99;
mem[416] = 144'hfbcee52fdc82022cfe4bfb3ffb90fcbdd868;
mem[417] = 144'h06eefe56f75dfe570d62f8cd0d9afdbe0048;
mem[418] = 144'hf224fdb2fb37fff70cddf0b3f457f20cfc21;
mem[419] = 144'h0b9ff541f0eefdd204fbf9d3000dfc82ef01;
mem[420] = 144'hf7aef5abfd450843ffe108d1055af2fc077d;
mem[421] = 144'h0c60f4710883f142f6f9f2bd05f2fef3f524;
mem[422] = 144'h0388084c065cfbc401a303db022efe61fb0e;
mem[423] = 144'hfbd8f283efe00718f89d0611042bfe1cefc2;
mem[424] = 144'hf524f953ee980c890228fe6bf462f9cdf467;
mem[425] = 144'hfe1df301fb1bf905f31cf351fde9faa3f87b;
mem[426] = 144'h0099042001290d7bfd34ecf4ee53f77d0422;
mem[427] = 144'h081b016206330d8f02610a3ff300fc340601;
mem[428] = 144'h00e6098eefd8f2eaf74cfee00924061309bc;
mem[429] = 144'hf448019d07e806fbf7b8fd2c0ed1070800c6;
mem[430] = 144'hfb51fe95ee0ef147056507e5f314f732e0a0;
mem[431] = 144'hf83cffd3efa9fab70947032f0149077bfee7;
mem[432] = 144'h096ff87c06650a7408dbf9a303070e3c0278;
mem[433] = 144'hf97d011bf2b1045e0b05f1cefdd30f9af482;
mem[434] = 144'hfb8ef74b0c19ffcdf9950838f96303840d47;
mem[435] = 144'hf04604e30a0b05d90d3ef1b9033704c5f563;
mem[436] = 144'h011e0c100076f97504bf000bf47f09c8f641;
mem[437] = 144'h0522f019fae0f72b0793f448033f011ef84b;
mem[438] = 144'hf8e806810908066deff9f0e10f9d055bf0fa;
mem[439] = 144'h00510a7f077b0278f689f541f8320bfe0461;
mem[440] = 144'hf7fff72af643fccbf43df1760964041d09c3;
mem[441] = 144'hfc5ef7fd00fe0ba9f88cfbfef1390a870ae3;
mem[442] = 144'hf5160c2c0680faccf3b1083f08c401d10303;
mem[443] = 144'hf18af01bf239fd370563f0370145feb40753;
mem[444] = 144'h09a50491f9c4023cf1a6ff3a09710ebff04f;
mem[445] = 144'h0b790894f6b40dc5042202bafd760625fe93;
mem[446] = 144'hf59903420765ff770a91f03f01e00453fd38;
mem[447] = 144'h051bf427f8ebf9f904dbf513fd45f72f0475;
mem[448] = 144'hef1b0a820658023ef8220ebafa64f82e0933;
mem[449] = 144'h0956f14ffc1afc32f7b606180578065c09ad;
mem[450] = 144'hf6ce0810f4d409eb0b12f583097e07b9f0c7;
mem[451] = 144'h0273fc2a06b9fe62fddc02db0753f46fed54;
mem[452] = 144'hf1c5ee7cf3fbf2c403f0f96af7f4fc24ff09;
mem[453] = 144'h03e708eafeed0d3eeffc0dab05b9027c0e1f;
mem[454] = 144'hf43ffd40fc53fbfe09d4fbd4fae7fc560f61;
mem[455] = 144'hf81604ddef3a07eaf3ea0c04f023f21bf46a;
mem[456] = 144'h08ca075f06e20d1c0653056df80503150c1f;
mem[457] = 144'h0c9c0797f590f5d2fc8c0c82f87ef2470296;
mem[458] = 144'hf80efe7cf34f0a02017bf597efb0f0fef84e;
mem[459] = 144'h047407550b9b099a02c7f55ff190093a0024;
mem[460] = 144'hf6dffd280b9f0931f0fef22507aa010cf670;
mem[461] = 144'h0211005a03f10df0f41308b6f02ff831f122;
mem[462] = 144'hfb2107dce9f7fa1cf5d00b1e06d107d70b20;
mem[463] = 144'hfa2a0b1e048dfd35ee96013605faf64a0b95;
mem[464] = 144'hfb6906e008aff3d70dddf607f189f369f222;
mem[465] = 144'h0caefda8facaf14dfbda0430f04efc49f0a0;
mem[466] = 144'h0b0f050c007c015509ec003c0345f7e1fb49;
mem[467] = 144'hfff7f65dfd69015e0607fd560219f705f8c5;
mem[468] = 144'h045800b3034c0563fcbdf4ac07fd0be50605;
mem[469] = 144'hf713fe38fb41099cff76010ff8c10ac3003e;
mem[470] = 144'h00a8fb45098702b907dbf52100b1047ef303;
mem[471] = 144'hfc3cf17e00dd065bf16f07def6b90742f40e;
mem[472] = 144'hfd3701200b1cfc85f7be0948fbc9f0abf3ff;
mem[473] = 144'h0c67f4960887f1e10e6c0da3feee0facf321;
mem[474] = 144'hf5f300a0ec08f986095defab0805fa7d0261;
mem[475] = 144'hf649f6d8f6a00c780aa000b1f7840602f17a;
mem[476] = 144'hf02c037df715f43300940075f310f30bffec;
mem[477] = 144'hf29afff7ffc8f696f7f5fad60ed80ee5fc7c;
mem[478] = 144'h04fe0631f7fc02310657fcdbf38d06b2f1c5;
mem[479] = 144'h0e7f030ef8b2fc4bfe04f5d3f167ff62f4e6;
mem[480] = 144'h06d3054e0976efad0f36f2e70fedfd4f018c;
mem[481] = 144'h0835f6f00b1c03e407610499f4cc02d50aff;
mem[482] = 144'h03eef5050e3ef5770a9202f10518f87801ef;
mem[483] = 144'h0e5dfff5036d0684f8e4ffc4f89eff420b8e;
mem[484] = 144'hfecaf1e1fe45f6290025f27ff972fe13f19d;
mem[485] = 144'h0b8bffe3f2c80c84f4c4f2d806db00d90aa2;
mem[486] = 144'hf8290b82f1b7f9a7f316f966fb3a0eda0a58;
mem[487] = 144'h08f5f617f769f977f521fa8f037a0a9efd98;
mem[488] = 144'hf90af8c00be00e0f0299fed6f071f12dfbe6;
mem[489] = 144'hf37cf8d306b104800915069efd60078e087c;
mem[490] = 144'h0682fda50919f27402c2f619f7d6fbacf580;
mem[491] = 144'hfbe8021bf78efddef71bf971f2090d25f247;
mem[492] = 144'h0dd90afb07f308df06b4fd530ae3075804a5;
mem[493] = 144'hffb90c84ff3efd89f83d003a0c8cf8190bd5;
mem[494] = 144'hf19ef6e2062ef4af0b3bf6a4f6f5f0dafdc2;
mem[495] = 144'hffebf21308090b4a02340db0fb19f83ffb00;
mem[496] = 144'hf45c0a99f793f686f2af0632044201830d9f;
mem[497] = 144'hfab00d610f7af6d109050c3d0cc70256f770;
mem[498] = 144'h0768f48404e8f424fde5f7a003b6feea0835;
mem[499] = 144'h06240d10f9850c1ff84f0e0efe240d6f0ae9;
mem[500] = 144'hfdfaf948ffa0f5f6f74cfecd0446fd28fd76;
mem[501] = 144'h08d6f72b093e05590a410a710cb30f20fa5a;
mem[502] = 144'hf28b07e5f5d407470c80056cf06cf5740e12;
mem[503] = 144'hf335075afe0d00080acc0c7df846f2ddf696;
mem[504] = 144'h0c3df2e40e39fe81f181fcbb0301f8dc04b4;
mem[505] = 144'hf0d3f14c0b13f1990368ff93f6920e97f7e0;
mem[506] = 144'hf58df469fff0fb62034f0d660e25f8c307bf;
mem[507] = 144'h0b49fcd205d9f47ff675f8a103a901150025;
mem[508] = 144'hfc53f79c0518058af6b60ebb02130a26f5e6;
mem[509] = 144'h0f15f83108e40071f5120ddb0e19ff03f61a;
mem[510] = 144'h0fd9fc3cfc66f3e4f219ff7109e3f6d800f6;
mem[511] = 144'hfb45f2580d59f02a02e502a60e3df4b6fa46;
mem[512] = 144'h034afd14094cfe34f9e2f2d6f737f0bff5b5;
mem[513] = 144'h06df05fef18403bff057f539f169002507e0;
mem[514] = 144'hf4cb04dbf0ae04970143ff87f84bfb6b06e0;
mem[515] = 144'hfe59069bf0be0b48fa51f2f3fd86043708eb;
mem[516] = 144'h08b3ff2afe02fae00126f24f070a0285f1a0;
mem[517] = 144'hf3f2f4d9f6e207820786ff2ef130fc03f68e;
mem[518] = 144'hf16bf930f889fac1fb490c24fdcef3e10a7e;
mem[519] = 144'hf4c1f4d50939068df9b10a8afac6f9ff0992;
mem[520] = 144'h0b800062090df1b2f2cd02e7009ef223fec8;
mem[521] = 144'h054c050afc90049b0297fb350a820f58fe00;
mem[522] = 144'h0224f68ced4f0569041bff860257f999f098;
mem[523] = 144'hf8bef43f015c0745fd4afa41f2550855f2ef;
mem[524] = 144'h02e6f45bff10fd090113f620f7cb0d7c0404;
mem[525] = 144'hf1260b2f0d7d0163065bf2f3f9650cff04ae;
mem[526] = 144'hf902f18807d7037d02d1f23afada08d2f66b;
mem[527] = 144'h05520b680c6f0c6bf7f402640d87f7c500b7;
mem[528] = 144'hed13f436f0e4ded9ef97f614e8bbf919eace;
mem[529] = 144'hf0b2f263fab1fbb4f6a704cff09ef35ff0b0;
mem[530] = 144'h0d2a0227fa1ff4c10b7c0cf20b71fe0dfac4;
mem[531] = 144'hf719f261de8dee6dfb8efb6af8a4feeef980;
mem[532] = 144'hf091f0fa0476050cffd700fc0399fa39fd64;
mem[533] = 144'hf6fe0baafc440b5ef3a80c39f989f88704e4;
mem[534] = 144'hf217f7c20d120e93f3f2f1acf7bc0ce0f487;
mem[535] = 144'hf0c7f7b60850fffb05def532fe4af475070e;
mem[536] = 144'h0829f71e09d201aff4f20269ef0d0106f038;
mem[537] = 144'hf3f6ffe702c4031902710cbe09dffb06f93a;
mem[538] = 144'hee6f02ebfdebfb920773efb9f3e1f643f62b;
mem[539] = 144'h002e05bff565073506d509d5000d07d709a3;
mem[540] = 144'hfe43f265f4a6fb8ffd4c032a0d61f92afa27;
mem[541] = 144'h0ad20213f99c01fb0d21015600360228073a;
mem[542] = 144'h032501d0e1e1f646e8dcebc0f522f59ce841;
mem[543] = 144'h0281f244fc44f03aef1c0463fc0d07fa0437;
mem[544] = 144'h0794fd12f1d608eff4aa02e5f52e09cef0ac;
mem[545] = 144'h0245faf70e1d0818f037fbac0068f8890510;
mem[546] = 144'hfbef03390956fd090213fb69ee33fd0f0bad;
mem[547] = 144'hfa32090b0153f7eefa0a05eb0a9f0a0e020c;
mem[548] = 144'h02fefd2ffa1ef98c05dd093a02d7eff1ffc1;
mem[549] = 144'hfec90c8df6c3f4950905f3b5f55afd15f27c;
mem[550] = 144'hfeb7fe88f4e4fba9085ef3dc0495055df548;
mem[551] = 144'hfd520ac10d9a04d70c580716f8600937fe0e;
mem[552] = 144'hf00106d5f36df620ff81f25ffa55f7c7044e;
mem[553] = 144'hfcc9005bfd79033a0988022efc47f7a7ef7f;
mem[554] = 144'hff55f4cf04e903a2f623029cfc65ee8dfec4;
mem[555] = 144'hfac508470be60911f39cf8d5fddf056e0620;
mem[556] = 144'hf6750217eef8005b0963039402d6089a0bc2;
mem[557] = 144'h090503010433f2d0faad0bcd0beb054c07aa;
mem[558] = 144'h088d0b9804f5ef8a0ad9f6e90a91ef2c01e4;
mem[559] = 144'h0da5f59cf56f099cf40507f4f020f11b0812;
mem[560] = 144'hfcdffaaef40804510135065b0365f224ffac;
mem[561] = 144'hf143f7f0fcad0a6005030562f96bff7df4ae;
mem[562] = 144'h0195f23df8f5055bef54f174fa1bf59bf3c0;
mem[563] = 144'hf7e4051ef90e03ed0402f453f3a0fc41ef10;
mem[564] = 144'heeef02450553f74a06cfefb8f842fabbf445;
mem[565] = 144'hfe22fff8f25a05d8f7cdfcc4ef9805230094;
mem[566] = 144'h0114f532fa0dfdd2ffdf0117fc8e03c2fa61;
mem[567] = 144'h0d86060efd800263feadfefcfa9afdb90bf5;
mem[568] = 144'h035aee280c9106f1fe9c0779f9860006f758;
mem[569] = 144'h05a701aef75601100ca4f7eef67e078bf1ae;
mem[570] = 144'hf0c5fd96f90d0c30fd7aebc0fd12f2ac120f;
mem[571] = 144'h0d21f092f32906d003c2ef65f35700d40d16;
mem[572] = 144'h04fbf32cfcd807000897009705f2fa3fe493;
mem[573] = 144'hfa5c00f0f2e7077af28f014efae702420e9d;
mem[574] = 144'hf09fea4cf19beac5ed4cf4c50214e71bf692;
mem[575] = 144'h0c14ff77034cf7740a30ef60f7250156fdd1;
mem[576] = 144'hfe23fc34f5c9f725fb3f0c45f5dcf2f6efd1;
mem[577] = 144'hf16ff904fb6808500bb4f932f6bcf3f50f74;
mem[578] = 144'h094f096e06be04c1f8aa035d02abf43b0c51;
mem[579] = 144'hf2affd3bef160b550789efd7fff3fa910610;
mem[580] = 144'h01fe06b2f4a50495f5f7fbd106c70b9b0a9c;
mem[581] = 144'h0ec1038401eaf5cd065f05e4fd56018404f7;
mem[582] = 144'h0b64fea6fa390393f8f10cab0cd709f30512;
mem[583] = 144'hf2fbff1bf772072cfd05fc24fce506010817;
mem[584] = 144'h0a6d0098fc7602e3feaf08fcf32aef62047d;
mem[585] = 144'h004e0590f6b4f5ed0c4402acf37bff1bf18b;
mem[586] = 144'heedceb34fb66071bf5fcfcca0257f8400e95;
mem[587] = 144'hfb29f722fa35f5c5005df437f93409bf0061;
mem[588] = 144'h082004b3f160006c03ca08d80aa7f997f8bd;
mem[589] = 144'h082e0b5ff4b405d702f8ffb0f51105900a0a;
mem[590] = 144'h0b3bed41f32af34809f2f2fd0a97067dfbf2;
mem[591] = 144'h0803000503dc0992fa130c3ef09def3efee0;
mem[592] = 144'hfad20a59fefbfce4f3bc02bffcce0567f552;
mem[593] = 144'hf13601dff30d05ebf898049c0c47fcd5fff8;
mem[594] = 144'h05650369078af93af41df5790ce7f85df7e1;
mem[595] = 144'hfe57f813ff84efd2f741eeabf55604cdf036;
mem[596] = 144'hfaee0ec7fef8f984059b006d07e6feda0687;
mem[597] = 144'h0809033aef86060cff3b0bb2f15f04dc0d5a;
mem[598] = 144'hf8f30d560a0a086ffce0eff9fce002f30d82;
mem[599] = 144'h099ef1a5eff903e1f699f2b50e19ff7500e8;
mem[600] = 144'hf7cd0510f4a6f351f3e7f0a60003f189099e;
mem[601] = 144'h0112f9cd098e0914f511015ffe670addf319;
mem[602] = 144'h01a1f59ffac5f9150aef016303a90269fe79;
mem[603] = 144'hf679041c0a580698f71bf8eaf512f7db0bdc;
mem[604] = 144'hfa72fc19f62af2bd0a9b0a05f08909fcfa4e;
mem[605] = 144'h0b47fab30ae80984f36c0e16fe34f148fbc3;
mem[606] = 144'h05a10b30f9a703eafae8ff8bff6c0152f872;
mem[607] = 144'h0b67fc9ef642f2f1f6c3f269fb9e02180ee2;
mem[608] = 144'h0e54f007010eefd2f5100b970cfa05f10f03;
mem[609] = 144'hf0d1097802dafd75062afb8105db02f90138;
mem[610] = 144'heffe0dc5f742089506a50432fea5fb1dfd31;
mem[611] = 144'h08bbfa4dfa3bfa40f506ef75ffe4fdd5f4b4;
mem[612] = 144'hfb7bfcc6f63b0e530c07049605a0f53a051c;
mem[613] = 144'hf7bef946f78b076107affee40ce5f4390943;
mem[614] = 144'hf02000b9f4f2f84f076dffcdfd6bf925f4f2;
mem[615] = 144'h0417ff21fff5012efbf6f5de02fff95ef6c3;
mem[616] = 144'hf23e083df4c2f2dffa56080f0c5607f90377;
mem[617] = 144'h08400be9f350f291f52700020e83f91ffbb6;
mem[618] = 144'h0cd5f2abf33dfd6a092b0954f09005c4f81b;
mem[619] = 144'hf8d50698fa780203f950fbc60e14fef20be8;
mem[620] = 144'h048e0b0dff7cf05efe88045ef28e05e8f509;
mem[621] = 144'h02c6f1bff47508f40073068ff86ff4d90661;
mem[622] = 144'hf0340e2701b203ff0778ffc1febff0020e13;
mem[623] = 144'h0f8df24607840228fe300d64fec9f87cfd2e;
mem[624] = 144'hefad0ef7f540f8fa0c190547f59cfc620227;
mem[625] = 144'h0deffe57f3ee0403f4410cfafb3f08e0f7f5;
mem[626] = 144'hff6404810cd0fb50f129fb3dfcd9f71cef55;
mem[627] = 144'hfe78f6ebee69ed370a7df8b0f4b8049d0425;
mem[628] = 144'h063b0adef4caf323f806f329f546f53b0e38;
mem[629] = 144'hf2190b9b0eb8fd37f5b8f269fdcd0e82f390;
mem[630] = 144'h010f02310025f549fbadfe7bf464f1010d30;
mem[631] = 144'hfef3028df6c602810f15f12efdb102cf0068;
mem[632] = 144'h0298fc80ffd9049ff0b2fbc40e8af094f0d7;
mem[633] = 144'h0af0efbef243f4cdf072fe6b07dbf483ef78;
mem[634] = 144'hff5cf99f07b5fa86fb130937f672f361f9e9;
mem[635] = 144'h0623f82bfdd8fb000975f6200a10f9c000ad;
mem[636] = 144'h041e080e0975fe19f95c00490a060c89fece;
mem[637] = 144'h03e8f8d80df20168f239f7520eedf0c90931;
mem[638] = 144'h0f4002b002caf213065bf3c50111f3ec068c;
mem[639] = 144'h0a16fe89fc81fedcfdf50d1002e8efcffa6f;
mem[640] = 144'hfc2ef6e0f911fef50d7208f8fe35f4f90a23;
mem[641] = 144'h0079090dfbcaf25ffbc4fc4ffcacfed7fbf8;
mem[642] = 144'h0f66f7bef573f2e0fdf7061b04c8f033015a;
mem[643] = 144'hf9dcf63b02e3fb0809b6f56b0077f220f9b6;
mem[644] = 144'h060af59604e40ca70aa807eef995009d0bd0;
mem[645] = 144'h0974f00607690b090964057800b40a4407a9;
mem[646] = 144'h03b50b8dfbf80efefa670b44ffe80b6709aa;
mem[647] = 144'hfeaaff53fd710938f8c9fe46f89803def33d;
mem[648] = 144'hf0e3f797f5b5fd67f1d7fd030738001d01a6;
mem[649] = 144'h0d0e0a170407020bfa8a003b0f9df0330797;
mem[650] = 144'hfc84079d08edf8ebfa66fcf3efb00817ed4e;
mem[651] = 144'hfe20f81a03730cc9fc000d6f044effd2fdb0;
mem[652] = 144'hf2c90f91f3770b7ff6cb02e80506f35dfd65;
mem[653] = 144'hf548fc93fb79ff3c0a64f214fa8d0a6207ba;
mem[654] = 144'hf88dfc85eedff9c1008c08e309be05ba04fa;
mem[655] = 144'h0df0fb25f95b0175f6daf7d9fb15fc3af511;
mem[656] = 144'hfd98e582f626eb51003501050126ff1ef761;
mem[657] = 144'h07cbfc900d89fb8c0a450592f6210471ff12;
mem[658] = 144'hef65f021093f065304c5f15207eefd37f991;
mem[659] = 144'hfa93f627f7cdf839ed7bf64f04e2ffd4fc91;
mem[660] = 144'h0756019c07a80bd907f0fbabf7e809ac0bc3;
mem[661] = 144'h0509f353f0d607790a7af2410dafeea1fb53;
mem[662] = 144'hfbccfd5f0d040915f4bc0410fc3cf19af516;
mem[663] = 144'h00690951ee7c02e0f3150ce407c9077b0ca6;
mem[664] = 144'h0053f26df7e6f4b6f0bbfb10001df25d0b70;
mem[665] = 144'hffa002c40809f7b30633fe76f05e02e3fd45;
mem[666] = 144'hec72f074078a011ceb7eff80e9dcf1fff49e;
mem[667] = 144'h06e3f9adfa9af641f9b70e0b055f0b70fb03;
mem[668] = 144'hf861089b001109760294f854039203c1fe5f;
mem[669] = 144'h02190ec20667fc240f4d03db0e740519f922;
mem[670] = 144'h0988fa8bfe4bf303fbce0465f75cf28ffac5;
mem[671] = 144'hfa1ef400ed6b0cdeef78fccb07c000a20205;
mem[672] = 144'h039af3dc0a2604e5f04df00202bd0a8c030a;
mem[673] = 144'h02bc076705dafdd5061507f6f78507e10013;
mem[674] = 144'hf134f0d2fc9606ab0181fa6dfc0d0cbc046a;
mem[675] = 144'h0619f788fac2f1c605ed01b8f900f6fd07e9;
mem[676] = 144'h022bfe5f0282ef33fac5f0da0f67efd805d6;
mem[677] = 144'h0d32007bf0d9f543f47df1b10904f0f8fa60;
mem[678] = 144'hfed8fa1e0e28fa04fbb8f9d5f989ff4a022e;
mem[679] = 144'hfb7ff11d0295f0baffa500f2fca903ea07d9;
mem[680] = 144'hf6ecf9d6067dfc280198fa020fb80797f9d5;
mem[681] = 144'h0bb30f450e18f8cbf0a101e100d00598f708;
mem[682] = 144'h0500efd1074d0b84ee470369faabfbb8034d;
mem[683] = 144'hf276fe9406de0c87ff9b0bd50422009b0e2d;
mem[684] = 144'hf3db0cc10148f16f05520b2ff8f5f6390008;
mem[685] = 144'hf42ff3f3fe2807cafbb7f79205280155fd84;
mem[686] = 144'h0637fae4edf208b2f946f3e7f3fefadffba7;
mem[687] = 144'h008e04fd079b0b54ffb501a70f320c6c06f1;
mem[688] = 144'hf232ff3c02e60d0dfd54f65b0545f47300e7;
mem[689] = 144'h07a5fb70f7c6fd05063cf6610c4cf5d3ff01;
mem[690] = 144'hf34f06fc08a6f295f5b0039cfe8705040dd4;
mem[691] = 144'h0cb10f5b0978fcbbf42401bb02eff726f764;
mem[692] = 144'hfe8dff01f846f110076af1f70923f539f2a1;
mem[693] = 144'hfce0f357095efdb4063f0f9b00c6f2ab0cc2;
mem[694] = 144'h0a2b082a0fcffaa502dbf1d808e20447f229;
mem[695] = 144'h05dbf9b0f8bffaf30777f0d6fb9b063ffdb1;
mem[696] = 144'h059afcc00eb9f9e30109fe63fb10030f0a4d;
mem[697] = 144'hf47df9180caef91cfb23052dff310fb8053d;
mem[698] = 144'hfbe9f0710896f689ff9409c2f048f46ffce4;
mem[699] = 144'h0aedf88b0cfb02c902e1053ef301fc50ffea;
mem[700] = 144'h09a1ff710c3808b0f0c7f7ea0cbb08edfad3;
mem[701] = 144'h0bc907590479f0cc00ebff6c0d23f2200833;
mem[702] = 144'h09e10c16f533f8e3047afd01082e06fafedd;
mem[703] = 144'hfc05f4d70bee012e07ffffb90ca8f1cdfc53;
mem[704] = 144'hf4900c0a01b80217f3e8fe05f8870d13f524;
mem[705] = 144'hfa380e4107b0f8bd0b4d05b40d7803b7f4ec;
mem[706] = 144'h034ff7b1fad50789f2b30f73049af48702ce;
mem[707] = 144'h0809ff63f3e6f10d02bbf6df0adef7870a3f;
mem[708] = 144'hf60afbc9026300c80204f051064ef485f7d7;
mem[709] = 144'hf81df0e2ef98f22903def775fa19f9b5fe0d;
mem[710] = 144'hf2a90ad8fc04f691faf2f3f7f3fd06f50f0b;
mem[711] = 144'h0de6f0260ca8007ff9ee0400fd46f5060030;
mem[712] = 144'hf097fa9403e1fa9c02b2f042fbac0c78f23b;
mem[713] = 144'hf84f02160279faf908a5fece0e6709c60784;
mem[714] = 144'h01eafa4efbef0344f0c70221f8bdf2f3f6c0;
mem[715] = 144'hf922029a0eecff9df5e5f099f44d0ee3ff1b;
mem[716] = 144'h0585ff340fac0ac704ec02f401e70190fb69;
mem[717] = 144'hf8e30f4c0624f85e00e2f167f40cfd1c0761;
mem[718] = 144'hf8ea0e66f204ffd3f9ec05fbf3b6fc77f1a2;
mem[719] = 144'h04090d51f2f3f2e100740546f3d8f1edf071;
mem[720] = 144'h0451f8de076ff82f0e5601d4fcdeefe9ffb2;
mem[721] = 144'h0b1a07f2fa6df763f967094f090208a1f6d5;
mem[722] = 144'hf169f47c0c71f2abf5fafe8c077af839f848;
mem[723] = 144'hf3ee04270608017807c8fc1e0c7d0dad0cff;
mem[724] = 144'hf506f47cfee50750fa1e02540a9aff5cfab2;
mem[725] = 144'h077df9bdf660f519efe809fe0aa4f4ccf4f6;
mem[726] = 144'hf2240264fbef0588f8ab0e210137fb2af751;
mem[727] = 144'hff9b0a1f0b12fa6ef1e404dd014e0e9af867;
mem[728] = 144'h0afdf7eef66f005ef7c4fca2f0400a1201d2;
mem[729] = 144'h062ff1f80401f676ff67fbe1045df949f647;
mem[730] = 144'hf4ea0386fcc8ffca07f5f08b0a02fbf3fc5d;
mem[731] = 144'hf0220c4f0b35fc8d0644f8dafa22efe80ade;
mem[732] = 144'hf5fefb76f0dd07e20bfcf9600f64f6050522;
mem[733] = 144'hf59f0389f69608caf75b0c02fa13057a020b;
mem[734] = 144'hf29409fcfdc8fb89f25eff5b084107c6fe3e;
mem[735] = 144'h0fd80360f8adfd4afacd065bfe5cf729ff4b;
mem[736] = 144'hf6d208d6fb950d12f84cfc1f0992fdf00189;
mem[737] = 144'hff9cf05afba7075904b5070ff7acfd30047a;
mem[738] = 144'hfd54f1230b440c7afbcaf816043c09000c9b;
mem[739] = 144'hf381f45efeedf9bbf5e4fa2208c808c4fdd3;
mem[740] = 144'h0bde09b30b3f05bdfa0d0823fb85fbe40c3c;
mem[741] = 144'hfcc90cf9f83f021bff68f461f1e3f155fa85;
mem[742] = 144'h0a0a05110514f606f7bf0bc80b3e069c0c0b;
mem[743] = 144'h02540d14fd5002010b5402d3077304daefa9;
mem[744] = 144'hf6b00273f3dcf6ef07af002ff00105150dee;
mem[745] = 144'h0fa7f9ccf769f9baf2b7f5280d09fba5f3b9;
mem[746] = 144'hfff40a04f43dff5bf37808610273f8610ba0;
mem[747] = 144'h07fa0c020c7604cf0d7cf0e9f714f76b03b1;
mem[748] = 144'hf1cb0d23fd20fd070d44f8f5fed0f3710ea6;
mem[749] = 144'hfd73f66bf49cf85f0d60078d07850dbbf858;
mem[750] = 144'hf0a0095dfb2006daf16d03c60d41f7b3f615;
mem[751] = 144'h01a608b3074bf5070d2b0cdcf088f373f125;
mem[752] = 144'hf3c8f545fe72f2080c9804b00dbff03e0a81;
mem[753] = 144'hf3ac082affc40c24f98ef59b02acfe0c0365;
mem[754] = 144'hfb6209e0f4370c6a0dcaf130090d0746f08d;
mem[755] = 144'hf30dfe2efd6ef2b8f10007daf6ff0695fa6d;
mem[756] = 144'hfdb1f38705a0017bfcb4f2c80a8c08ac0700;
mem[757] = 144'h0140068d0683fa76fd400937f6910f69f19b;
mem[758] = 144'hf808fe93f407f8df0b6afd7afbdc00f804d1;
mem[759] = 144'hf9670e4cf6fbf774051400360f54f7890a3a;
mem[760] = 144'h086804caf12c0fdd08c40a6cf6ab03e30001;
mem[761] = 144'hf127f1e9fec6f6a7f3400d7dfba2fa300fc3;
mem[762] = 144'hf5620908f338f82dfb06f69ef17101cef2c5;
mem[763] = 144'hfa79f96cf214f7df0c080ffe0bc6f5230f95;
mem[764] = 144'h0c4ef1ebfc16f66f087cf308095201b7fd39;
mem[765] = 144'h018dfe33fc9af15af6de0b510c86fb6c060e;
mem[766] = 144'hf67202b7fbaf079cfe2709430f30f89a01f7;
mem[767] = 144'hf157f217fa670bb7f244003d0f3df25afec5;
mem[768] = 144'hf0dd060aff38039c0c1a02a5fd4ef642f656;
mem[769] = 144'h09fa0d1bf630089d0e34f349f630ff7af5b1;
mem[770] = 144'h06520ae205d3023206330212f0e30a32f70a;
mem[771] = 144'hf7e9f2c602ff05ad0798fa29031c0c88f2ee;
mem[772] = 144'hfc2208d70255f9b8f266f1cc078cf3e6f828;
mem[773] = 144'hf438034d087f093bf11a0103f82f0529f244;
mem[774] = 144'hf758f3acfd27041200cdf125fb28f5d1fc9a;
mem[775] = 144'h04ccf9e800d1f468f3f4f20d0757f61508b4;
mem[776] = 144'hf78ffec2faa4f14f00f3f79f07a80e88fa62;
mem[777] = 144'hf2e0f69efa3efbf20625f6280f92f594f552;
mem[778] = 144'hf944ec710a7e0287f4d40b8b01980c6ffdde;
mem[779] = 144'hf006f62e0974fa120a5506f8f680ff87f3ae;
mem[780] = 144'hf2930eeafb67fb7df6d8f6bffab502520bd4;
mem[781] = 144'h0b94f1aef0bdfbddfc12f044033bfe20f69b;
mem[782] = 144'hfa35f618fd9def0802b70da4013cf1bbf51a;
mem[783] = 144'h0858f4c7fc090d12f0f3f9190513f4430632;
mem[784] = 144'hf4f3f6720bdc0df208a3085bf956049700ac;
mem[785] = 144'h0512fb05f90cf10508f50a18f3d8f6d00ba4;
mem[786] = 144'hfb61f748f4c30b12f540f175f2f40dbf06c3;
mem[787] = 144'hf115fba60dd40625f045fd0c065b04d90835;
mem[788] = 144'hff56096c0bb6022df847046f04440503f3f4;
mem[789] = 144'h0e71f1df044306ee01c9f77e06fa05c9f47b;
mem[790] = 144'hfbadff12f3c1f2f104ab08de0eccf396fd0d;
mem[791] = 144'h0c4c088c052b0794041bf47d0eeb0ead0666;
mem[792] = 144'hf1fdf915f554fad20a7bf018090701dbffb4;
mem[793] = 144'hf0c403f909f302d8f2a9f89e0357fa32f68d;
mem[794] = 144'h0e4700e9fb690062f85ef078f2b70a26ef68;
mem[795] = 144'hf4d70bb7f57502b4f55dfcf9f70d088eef76;
mem[796] = 144'hf912fbe70251fab10fa60e6bf6caf87bf804;
mem[797] = 144'hfde003dff729015c08810723f54107d70afd;
mem[798] = 144'hfd85f602fbbb01f8f015099bf86a0150fafa;
mem[799] = 144'hf40e0cc0004e07c9f15e0131f3d40b1603b0;
mem[800] = 144'hf68fe68af511f62c05f4f56cf226f75bfc4f;
mem[801] = 144'hfc15f127f7bf007b0a240f3e05a3084e0021;
mem[802] = 144'hfa2906cdfb94f28306df0d47f111f438f170;
mem[803] = 144'hf293f622f971df3cfb65fb81ed4fe97dfc3a;
mem[804] = 144'hfe41f40106bd0ba8edc00b88ee46007f0769;
mem[805] = 144'h0168f517fb11edd00aeffc1f011ef58f01da;
mem[806] = 144'hf05a012bffc5f1e7f752f9cff9ea0491f457;
mem[807] = 144'h091503b10513f27cf3e60b11f44f0692ee9a;
mem[808] = 144'hfd23018aed1cf68df61bf7abfa44fcc5ff8b;
mem[809] = 144'h060107dbfb09023a0385f73af54ff652ffe2;
mem[810] = 144'hfbc51bd8efe9dcc5094805a7fe45125f0779;
mem[811] = 144'h0c1601490ad405fcf658fc9001e9fa42028e;
mem[812] = 144'h0a3af32df9e406e7f3e3eca60211064409ca;
mem[813] = 144'hf446066cf18c0abf045406f8fca60486ff91;
mem[814] = 144'h006bee35e39ff9b6eaa2ed23fea9f8f9fd6f;
mem[815] = 144'hf5650333f842f629f51609e1f5dc07b7f159;
mem[816] = 144'h0a5809b6027d0d3aef47ffc1f886f67cf970;
mem[817] = 144'h06840b21fd5f025e075c07d90c8effb00eec;
mem[818] = 144'h0548f88400ecf5effd17fe7cf49500730689;
mem[819] = 144'h0dbb089d0d4ef74af796ffc0020bfdb3027a;
mem[820] = 144'hfc4ef1da02210af2039afc420f0108940813;
mem[821] = 144'hf300f89406eb07000cf6f4b102c20740061e;
mem[822] = 144'hfc21003e0ca507530c2903eaf6f4f3b9f069;
mem[823] = 144'hefeb03b6fa65fce50b3bff07f65bfe150398;
mem[824] = 144'h026a0b210444fd43fc93f10ff142044f0c9a;
mem[825] = 144'h0330ffcdf8aff6acf4e50893f3470089f1f1;
mem[826] = 144'h037cfc3eeed0008ff5c8f2e80392056b0819;
mem[827] = 144'h04dbfa70fc9cfc36f12309c204e9f791f484;
mem[828] = 144'hf16f03480f39f1ac006ef13ff10603a10340;
mem[829] = 144'h00010f22fc150d0a09a40e0b0b62f9fcf259;
mem[830] = 144'hf18b05befaeb0bb0f27209fefe31f693ed5d;
mem[831] = 144'hfa47f7a1073e0917fcb20e1e0d74098ef851;
mem[832] = 144'h0840055efd9ff6450e3ffc23f84cf9e10036;
mem[833] = 144'hfd54f2deff13f7ba095a0d1307e1f30ff8ff;
mem[834] = 144'h029dfa98012df15e06700bbf0a9cf8c5f779;
mem[835] = 144'hf5120becff14f2d7fa86f0020d54fde9f5d2;
mem[836] = 144'h08d6012bf4fff93c0c2e0869082b0285f791;
mem[837] = 144'h0085fc5f01eef403003ffe0bf77c08ba07fc;
mem[838] = 144'h09c90176062bfa700eb406a20de508c1f250;
mem[839] = 144'h044cf42c04c6f8a10ea60327086a0480017e;
mem[840] = 144'h0ede0b84fef9faa5f3a0f21df5db0968f735;
mem[841] = 144'hf033f1d802c0f5c4090301e10fa4f027f9d5;
mem[842] = 144'hf18cf24e011907b6f1e00d4d082cf492f0db;
mem[843] = 144'hf6bcfb6901bcfb3cfbd0f64ef037f725fbc2;
mem[844] = 144'h09cbf94207f00a770f1b0df9fb1205a8f682;
mem[845] = 144'h0890082f06e2032e0034fc3a0b53f908fe39;
mem[846] = 144'h0a74fd9e042ffa06f407001ff3acfb18fb05;
mem[847] = 144'hfa090c790d39feecf7daf5090371010dfaf6;
mem[848] = 144'hf40f0e1700adfffef1fc0efaf401f1e00654;
mem[849] = 144'hf198013c0d96fc6afcd2034c09e9fb1f0e30;
mem[850] = 144'hf767fa47080005eefa8b0d860175fc45fd01;
mem[851] = 144'hfe01f3a903c2efabf51bf20af214fdddf8c3;
mem[852] = 144'hfce4095c0c90f7d0fb84ffdbf9c806210914;
mem[853] = 144'hf700f247068e014b0878fd49f4bdf42aff40;
mem[854] = 144'h08a9f91a00b1036afdaa0c5404f3f569f479;
mem[855] = 144'hf1ce0c86f554ef2d00acffe10db2f637ef28;
mem[856] = 144'h05640a1e095e09d805bbf2620225f3a103b2;
mem[857] = 144'hf3560a61f6af09e2f64a0e42f84bf454fed2;
mem[858] = 144'hff1902d8f2b80b0dfdb8fa3203befe0cf540;
mem[859] = 144'h03090c52f3d1f5e70757f6660e260db80c14;
mem[860] = 144'hf9520428f8dbfe18f6e5066e062c0d6cf68f;
mem[861] = 144'hfe1d081b06acf22af21f037704a90d44f2db;
mem[862] = 144'hfc5ef785f3d6f0370980f492fcf1fbb7f302;
mem[863] = 144'h01c3f04ff226056dfdebf0d801b0fd03fb9b;
mem[864] = 144'he5720403ded90303f6db0d9fe8afe414e022;
mem[865] = 144'h01f30cb308c40829f37afe26f5f709c301b7;
mem[866] = 144'hfb6cf13f05f6f8b00153057bf44ff63bf6f9;
mem[867] = 144'h02f5ef06f659eff1fd44f1d3f4090614e8e1;
mem[868] = 144'hf1d602bd020601e4f4caf71aefeb06affbbc;
mem[869] = 144'h08de04d801770d17ef66f903f5a5fa39ef66;
mem[870] = 144'hfbeafb98035ffe170b16fda1fc8600da0eb4;
mem[871] = 144'hfc6a0946f7010c51f75ef9bc09490d4b0e62;
mem[872] = 144'hfbf20730f034feb40b6a03090c11f17d0180;
mem[873] = 144'h0c5cfa58094a07a003d3fb5c09f901d6fb85;
mem[874] = 144'hf871064b1243002c015306d2fa1b065a161e;
mem[875] = 144'h0692f465faaef65208a90b4309080b57f856;
mem[876] = 144'hfe4503e5f115f097f178edd1f0b0f620f271;
mem[877] = 144'h0d91075b0601f07afcfa0f56fe9d05b4f353;
mem[878] = 144'h0495ef11f993ed27f13cea3b0280fb000753;
mem[879] = 144'hf932fc6f04c9ec440a8df447f0d708120c0c;
mem[880] = 144'h0321fedf090df5e1fcf50c34fe4507820404;
mem[881] = 144'hf8ab006cf917f943f4b2f146fb8ff3ae088b;
mem[882] = 144'hf5f2f2100cda07cd0fd9fb670d46fb03f46b;
mem[883] = 144'hfe51f9ddf4ee036bf1a70b100c7a00f7f2cc;
mem[884] = 144'h039ef76a0536f8830b30fb48fe2e02b40acc;
mem[885] = 144'h0c270927f847ef2ff31f0d80f1eefa6d01e5;
mem[886] = 144'h0a38fbcbf32807800af00e7dfcb20353f4e5;
mem[887] = 144'h0d30f677028ef23bfd5103a0f6cbf6fa0cf3;
mem[888] = 144'hf125ffc3fa28fa49f3d70530fb4c0ec0f704;
mem[889] = 144'hf8d1f541f11bf92dfc1ff111f787f0c601eb;
mem[890] = 144'hf48e09fdf2ffebf20653f0d10866035ff1de;
mem[891] = 144'h0e01f780049901a00c8df47bf41f0d620768;
mem[892] = 144'hf31b0d1a0e6305d1f1a4f251077dfd38f437;
mem[893] = 144'hfc1e07a701fcfd6ff9ccfd0cf1e4f1ca0bfc;
mem[894] = 144'hf09bf584077603ecfeacf90e0bfbfaf004ed;
mem[895] = 144'h0d8c06840779fc2408d00b5804b5f0bafc5b;
mem[896] = 144'hfea90bf804f409ad0ec6fe25f262fa28ef84;
mem[897] = 144'hfce9f1300e6aff720a130325fd1c0478f1d9;
mem[898] = 144'hf818ff28feb90118055209a200dff41df8bc;
mem[899] = 144'h00caf75f02b60cdbfc5cf660f5aff40bfb01;
mem[900] = 144'h0cebf77c080e034a0706fe870221f785085d;
mem[901] = 144'h01d204ecf24ffbf1eff1f7b60ab60860f97d;
mem[902] = 144'hff59f939f3f203d3f5140171ffa4061a06e9;
mem[903] = 144'hf0fff3bb03f9fd87ef01f0d001360e9c0675;
mem[904] = 144'h0430ef34fc040b68fd9ff98df78b09b8f519;
mem[905] = 144'h0ed2fb24f345f2a0fead03ce0a13019bfbfb;
mem[906] = 144'hf3350669082d043f0099036005a8ef1affc0;
mem[907] = 144'hfab603440bb6091cfe00f85af53d0710fac3;
mem[908] = 144'h066dfc5bf06a082f09540a4cfa24fdddfb9b;
mem[909] = 144'hf0b8f395f6170bb60c8b0ec204c302bf0f85;
mem[910] = 144'hf145f5b8f5f901cd0b7d0ce3f0fb0b90efd6;
mem[911] = 144'h0dd3fd99064eff7b06c503f400b2028b0833;
mem[912] = 144'hfea3fc8cf606f36f01fa07ff0d2e00170037;
mem[913] = 144'h028cfe0106ff08bbf0ec08fc0dc9078902d4;
mem[914] = 144'h0afefbb6fc89fa580c6702640a50ef58036b;
mem[915] = 144'h072c0598fd5c087e07510264f9360d6d0aee;
mem[916] = 144'hf588f814faeb0120f7eb064a0091f456f841;
mem[917] = 144'hfa1f0697fe55fd2909320fbf0ba1fada0896;
mem[918] = 144'hf791f022fd2cf984f08705eefa930b7cf6f9;
mem[919] = 144'h08d10914008c0571fbcaf19c03ab0a5105da;
mem[920] = 144'hf2c8fc02f94cff310f520d59f40506b4f13a;
mem[921] = 144'h06cff44df47bf2730129fecb03b30b78fc79;
mem[922] = 144'h0a7df776032503c2095802eafa0a022eeebd;
mem[923] = 144'h0961ffc7f479fe01f1f0fb7afdbcfe5bf324;
mem[924] = 144'hf6defc5afdce0e8300b1f770f911f5e2f00d;
mem[925] = 144'h040cf3e508b204ddfcb7f8fa0209f63f0626;
mem[926] = 144'hf377ee94088cffd1028a04ce0f7bfe01005a;
mem[927] = 144'hfcc9fb690484f6ebfbacf557007afaa4fd7f;
mem[928] = 144'hf9b90b91eee6fd7bf8660ceef4510d6f00e3;
mem[929] = 144'hf9f805c00b16fe4801470a1ef324061a0c5b;
mem[930] = 144'hfd8afd250daf0d5efb5105b4f9e4fc95f036;
mem[931] = 144'h0e5c0dfcf5a7f259f72cf1c40518023e0363;
mem[932] = 144'h08c80629f6c3f2bbfb61023cf797feabf5c5;
mem[933] = 144'h0f450680fe8ef11ff9fdf1b1058d00bd0b1a;
mem[934] = 144'h0884f72b063d0d3efca400450e8f0154f79f;
mem[935] = 144'h060e0c94fb84fb7900e40c710e740217ff3b;
mem[936] = 144'hf9cb0b8700ce0e1a0190f0280bcef51effd4;
mem[937] = 144'h088bf1640518042d049607bdf9c205ecf0c4;
mem[938] = 144'h0934065e09c5f451fa5d01edfaf2ef23f883;
mem[939] = 144'hf5c50b370bd1f97ff85cf4eef1feef36f41c;
mem[940] = 144'hf356f30f05cc0ef4f6c4f2faf28b07720a14;
mem[941] = 144'h03f9fac8fdd409560663f5a8f4b6f223084f;
mem[942] = 144'hf5f503be00c3f1860207f9030e900c2b0799;
mem[943] = 144'hfb74f0e1f239f6000ae3043b05c60595f9fe;
mem[944] = 144'hfa0ef02f081f0bdaf3f3fbcff4f4051eeff4;
mem[945] = 144'hf48df85a00b20a970a39f71900d3f35d0041;
mem[946] = 144'h04e103b8f2e30a63fdd702a3f74cf8f103f2;
mem[947] = 144'hfc5dfaf7fd51f1eefd09eff9f6c30862f9f6;
mem[948] = 144'hfc5207e4fa6efbfa0860fede09b7fc14fba9;
mem[949] = 144'h0598f025f716ff660cdc0b72f75ffcc7fd61;
mem[950] = 144'hfd52f5c406afff90fad4f1d30be70d4cffd1;
mem[951] = 144'hefdb05560cfe0c2b0c40fc310e6908a6f119;
mem[952] = 144'h033af054fe6406b80087f575ff3ff21604e8;
mem[953] = 144'hff990025f391fea0f61d0cacf08f0f560b61;
mem[954] = 144'hf983f8dd06fff1e3085df5c1f911f3bdf0fd;
mem[955] = 144'h02a5ff9e03d7078af07df5070c97f9ddf902;
mem[956] = 144'hf084fedbfe22f01d0ed7f5f4f66df82bfe7a;
mem[957] = 144'h0dde0297f87904adf1a1f5770e3201860197;
mem[958] = 144'hfa080bb1f424f4ed0ea6f31e064defabf379;
mem[959] = 144'h03d4f9eaf0cdfefe01b3f7ccf71405360e3c;
mem[960] = 144'h0c3ff39a01d10636f49cf3a3066dfed50c54;
mem[961] = 144'h0f400c64f19005840dde075303a40e9800cd;
mem[962] = 144'h007d04ac01a9009507690d1305f7f551f61a;
mem[963] = 144'h042efeae02c7fa810e74ff64fe2f016e0985;
mem[964] = 144'hff3efad50f09018a0a86f80c078bf1160903;
mem[965] = 144'hf4d801d801e8f2330d19025802f00e190f9e;
mem[966] = 144'hf0c507b002d2f2c90779f9f0ffeff15defcc;
mem[967] = 144'hfee6fa09f7c60312f7d7f3a4f5c3f84607b2;
mem[968] = 144'hfc7cf2d107cb0bc6087b0944fa61f217fa51;
mem[969] = 144'h0f3508f2f1a508dff9710a5003e3fabdf272;
mem[970] = 144'h0a280cbdf4bc0ceef274f79ef50ffe5df4d0;
mem[971] = 144'h0c29033efc84005cf11b00edf695f3f3f8d5;
mem[972] = 144'hf73b030005720734f544071ffbf60c32f5d3;
mem[973] = 144'hf23e03aefb54062cf28df8e90738fb150927;
mem[974] = 144'h06ce071603f306a10806fa0704d6f6abf406;
mem[975] = 144'hf5da0c57f780f6f2053802e30ab30f28f578;
mem[976] = 144'hfd5c06fe049fff56f8660072043e03f00a3d;
mem[977] = 144'hf346fe790e80f273feb7057ff816fd33096e;
mem[978] = 144'h0de80434f9eff3e10fbd0ca9ffcf0228fc59;
mem[979] = 144'hf05f07b7036509a30c830403ff72049df643;
mem[980] = 144'h0bb20d29f691f0d004ea043605b8f074f784;
mem[981] = 144'hf62e0533f76206410d3b02abf8ea057309de;
mem[982] = 144'hfb39092c081f09e6f3b6fad0f31d0e53f0f4;
mem[983] = 144'hf7b00b8af2350e89064d0908f869f6c0f65e;
mem[984] = 144'h0d72f580055c02340bdf0b12f9540809f470;
mem[985] = 144'hf6b9f7aaf3c70729f611fa640f21fd9202a3;
mem[986] = 144'h065400040cb6087cf39afdef0643f185f07c;
mem[987] = 144'h0ceefd40f3e1fe60fac8ef7b04ad0e440d27;
mem[988] = 144'hff6cfea2f46bf5e807cb0278fcf9fd5e0938;
mem[989] = 144'hfd3ef47f0bd1f293f3ddf33efaa4015ff275;
mem[990] = 144'h00680b3b09baff750a0c02130186068df6e5;
mem[991] = 144'h0926021d018104500c0dfd91fee3f5970591;
mem[992] = 144'h077af9c9fe5bff09fd4cfac5fa56ffda0207;
mem[993] = 144'hfa8df70f05110ef9f1ca0eb9f5fd01b10448;
mem[994] = 144'hfa6bf98a0c9ff141fe99fe71f8850697fe2d;
mem[995] = 144'h0b2f0338023703bceb4dfaa0fc1006b1094b;
mem[996] = 144'hfb350cecfafdfd90f603f08e08ce01ff05be;
mem[997] = 144'h0613eeb3f0a5f8b5fd09fc31fcf205d702e3;
mem[998] = 144'hfda1f9a201ee0bd60dd701f901cd0ae901d5;
mem[999] = 144'h02f200eff3930027ef5e0926017bf173fe4b;
mem[1000] = 144'h0e87031305b0faa0f1e0097505d0f825f300;
mem[1001] = 144'h0faef09afeecf754f021f8f0043507eef2b8;
mem[1002] = 144'hf259f0a4fa67f74afce1020a0a9df419fbaf;
mem[1003] = 144'h030d08e30d6ffebded6cf45709900a8fff93;
mem[1004] = 144'h06070ac0f7f3f8810abc0709efc6f449f746;
mem[1005] = 144'h0a40ff00f62007750f99f798f3cff48af6a8;
mem[1006] = 144'hfd5f0d2bf11ff3fdfec907e10e73f92b02e4;
mem[1007] = 144'h0702fe3809da05030ab703b20201fcee073d;
mem[1008] = 144'hf59ff9230603f1b2fc7c0b1df2d7f6b00779;
mem[1009] = 144'hf0e6f59ef200019400a7fd0ffcfff2d0fec8;
mem[1010] = 144'hfb1406dd03320507fa75f5c5f09405fe08a2;
mem[1011] = 144'h0bb7f5e20976f139fdc7fb0dff4cf5fdf6ec;
mem[1012] = 144'h04100205eff8efe0f5d8f177fa86f987f823;
mem[1013] = 144'h0142fedff74bfd43f563ff74f4c0f35e0794;
mem[1014] = 144'hffb3fc2cfc210401f648f715fc30f1570ba5;
mem[1015] = 144'h0401f5efef74f4180770f74affe9035ef6e7;
mem[1016] = 144'hff1bfdf0fe3c037403a30a55fc3804caf09f;
mem[1017] = 144'h084ef0c6f5fb0b820929f71a0a07fd95fb05;
mem[1018] = 144'hf4170175f87300a1fd05f7befbc4f314fd69;
mem[1019] = 144'h0355fa15059cf4eaf1f8018d089c0a7e0dfa;
mem[1020] = 144'hf83afcbef3df029afd2304440d49fc0df2f3;
mem[1021] = 144'hf498fb910b64fcbdfdb0f123fac9f327f7b4;
mem[1022] = 144'hf9e1f6eeff5500f00211005f0a59f2440484;
mem[1023] = 144'hf757f81ff08df23a031ef5910153f10e08f0;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule