`timescale 1ns/1ns

module wt_mem0 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h035cf13df617f51cfe9c05ec0b70089d0243;
mem[1] = 144'h020905c00dc9f4e609310dcafa5305cdf2f4;
mem[2] = 144'hfee2ee7ef3df05fcefcafcdef6f905ecfbdb;
mem[3] = 144'h0a13fbbb019ffbfdeee006e2022e00b70c08;
mem[4] = 144'hf6def11006f10748079dfb9a00a1f3b104fe;
mem[5] = 144'hf84af7f80bf6f2bef92a00c404fa07e4090d;
mem[6] = 144'hfbbb069af91c05f0fddffeef0d5cf2e807bb;
mem[7] = 144'h0ae0f61cf9fdf5e40a17fb81fcc108980c03;
mem[8] = 144'hfb22095af14b0daaef550dfd0728ff6d017d;
mem[9] = 144'hfb0704e5f19ff0e4fffbfe9d0017f1ab02b0;
mem[10] = 144'h0499fccc07f607520738fc600b870051f7f0;
mem[11] = 144'h0b4b01e8f724009e04c1f4cc00bb0a71ffe8;
mem[12] = 144'h03c50bec0e07f8ce07a40970039e05c001c9;
mem[13] = 144'h01f50aa4f58403c9f022ef6cfb9a03a0ef4b;
mem[14] = 144'hf2dc064df3f5eef70306f96ffb7ef40bf630;
mem[15] = 144'hfec20cf6f9bfff7efddefbb20257033f095b;
mem[16] = 144'h08530c6aefaf00a60480efe1f8ecf89bf1b9;
mem[17] = 144'hf24e0c0c045b06a20788f141fd3303c80f36;
mem[18] = 144'hf5dbf6e90f190bd0f0530d8a0df00f570d21;
mem[19] = 144'h06a5ed46f265fbe000b9f2b30be9f7e3f0f2;
mem[20] = 144'h065bfb9201ffeec6f967f6aaef0ffe85f928;
mem[21] = 144'hf79404eaf1010573feb4041bfca702e80af0;
mem[22] = 144'hf24900660c3eff8bfd6d0b1b074c035902bf;
mem[23] = 144'h099e0d4affddf8830684f3690757f4ecfc47;
mem[24] = 144'h0e260210f3b1fac6f7190dd80b0af6d50368;
mem[25] = 144'hf3aefed1ef3df64401080ea7f2ff07d104ca;
mem[26] = 144'h00dff760096ffdda01bb0a86fbb802270cfa;
mem[27] = 144'h037af57b0d0703ddf0a4f420f43cfd09fde1;
mem[28] = 144'hf30e07f9f98ffc09fd28f2c8f0dbfa37fff4;
mem[29] = 144'h0ac802b60ddbfc84081b034ff8ad0d3ff9ee;
mem[30] = 144'h03940617ef9c040efcdcfc03f921fa2f09c7;
mem[31] = 144'hff1efeb2faad0b2009810438f5b0f005072d;
mem[32] = 144'hfe2e006700cf09d503a40b13f4ccf2b1f35e;
mem[33] = 144'hf812fd2f0e56070dfbf5f98bf064fe66f6b6;
mem[34] = 144'h0a65fae9f24b038c032905b5ffe0f8a90682;
mem[35] = 144'hf361ffe200c707ddfba7099af5d8f010f0f5;
mem[36] = 144'hf1650d7a01d2f8620e7c0d90ff9701af07f4;
mem[37] = 144'hfc4d03cb035afaaf1025f5660801f4f50796;
mem[38] = 144'hf1c9efeb0535fdc8f1e8f8770248f442f15f;
mem[39] = 144'h054ff31e0164f4a4f57afc96f6b3ff3b03b2;
mem[40] = 144'hfe590beef6420cfe068202c5fdeafce5f81a;
mem[41] = 144'hf7fb0a40efe10916f6e4fc2ff3f802d7fea7;
mem[42] = 144'h09d0fedbf66afaa0075f0d7df0d10b13fb72;
mem[43] = 144'hf4b9006af225fa4008fc02f1041ff8a90600;
mem[44] = 144'h04b3eff40799fa7500f9060805b5f578056a;
mem[45] = 144'hf0890953fec2f9b600d8f6ba0ce00abd0a7f;
mem[46] = 144'hfb5ffdfd05a2f1f60c9df38ffddc0a28f857;
mem[47] = 144'hfa21f0b2029f0ab8fab3f0c00ef8054b0c48;
mem[48] = 144'hff140eff02b0fab407750c1c0c21f2910c6b;
mem[49] = 144'h06f8f1eefb180a9ff80e0ca607f3feb9f9d0;
mem[50] = 144'hfd9b0a13069bfea2027ef0c30bc90faaeff0;
mem[51] = 144'h06d80d1cf6e403a60644068cf8730d55078f;
mem[52] = 144'h0145f285f545076afaf8f28e0e37015ff864;
mem[53] = 144'hffebff54fde40130fd4001adf998fad9fede;
mem[54] = 144'h0b41f2600c4d049ff1880d4bf2bcf108f2aa;
mem[55] = 144'hfdeffb48053d095d0092f0ecf67a00040838;
mem[56] = 144'hfd4c052df751fe3407b20d830293fad5f334;
mem[57] = 144'hf54c03c9f8c9fd42ffc3faceff96f4b8f3ac;
mem[58] = 144'hf02ff94bf333ef3df4c9f89e04b5fe3a0d38;
mem[59] = 144'h09cbfb80f3c6078f0976faae020bef8a0cad;
mem[60] = 144'hfd610aa40ad30081024afe3c09e902a3ef68;
mem[61] = 144'hf038fe15f748fb94f02a0603fd9aef8403d0;
mem[62] = 144'h0752fd6df5eefccaf497efeb04af0a41f014;
mem[63] = 144'h042e0172f522f706f9e60d7bff63f31df671;
mem[64] = 144'hf843f69b0c17fb450285feefff8d0e130d15;
mem[65] = 144'heecd00160985074ff2c5efb0fcfefa40f8e6;
mem[66] = 144'h0e28f2ecfb5af519047f05260345fae6f668;
mem[67] = 144'h077bf42100540f9c05c7faedf9650ab50e11;
mem[68] = 144'hfdecf43e09b8f239fc710bce07660aacf83a;
mem[69] = 144'hffdcf39b09e80d6af906f0ec0c0bf35dff9b;
mem[70] = 144'h0418f2bc00fc0e9afceaf979f8d2fe5007de;
mem[71] = 144'hf7c90a02013103660b0b0ab10b930ed0f9c9;
mem[72] = 144'hf07cf1e50a7efbbbfb700be3fc1b0ed105cc;
mem[73] = 144'h021900a6f753f535f46ffa9204bb02e909ee;
mem[74] = 144'h09c40976f699f753f58f03f00400f9610765;
mem[75] = 144'h02e4030cf88ff9be0dff0545f5dbfb43ff82;
mem[76] = 144'hf3fefd05098b0663f87c0acdef83fe620c8b;
mem[77] = 144'hf06af592febc00440a55f2fdfd5206a102fe;
mem[78] = 144'h0c69f0daefcdf7b00b2cf05afcf2f7060645;
mem[79] = 144'h0001063ffbed04650557fdc70f11081801b6;
mem[80] = 144'hfa78fdf104420518fdc2efb8f8e908330367;
mem[81] = 144'hff72f1e8f3b3f32cf925047e057ffbf10d6f;
mem[82] = 144'h0fb1f0f0f980f0cb00f3fab9ff2cf083fc0e;
mem[83] = 144'h0b93f4cb0b1dfc26f92b0ba508b0f1b70d60;
mem[84] = 144'hf8f8f19e05f2f27efeb8075e0f52092cf235;
mem[85] = 144'hf7aefd5df332faf8f7e30c8906fd0df9f0ab;
mem[86] = 144'h0889068afa4f0abdf566f013feb6006af6ee;
mem[87] = 144'hfa8f0cc7054402f7fc4ff56a00930549f6df;
mem[88] = 144'hff6208c00fe5f5c6fb000090ffe908620a2a;
mem[89] = 144'hf0e10a0bf07f008b0f880835f320f6b404e0;
mem[90] = 144'hfe18f60203b30420f51df22e0e44044e00cd;
mem[91] = 144'h00d80b440779ff9dfc680c1e06dc075704b0;
mem[92] = 144'hfc5ef4e7f1c6010ffbc7081a0b6af2f5ff67;
mem[93] = 144'hf5fcf5b6f6e5f65f0804017d075408daf88b;
mem[94] = 144'hf50303a503d8f438fe4df884f257f2f400fc;
mem[95] = 144'h04b3f9d10c8af68b0d8b08e00d1502fd0669;
mem[96] = 144'h021a06d3f2e6018403a3019f002cf822037b;
mem[97] = 144'hfc57f22cf2650507f29807100587063af87f;
mem[98] = 144'hf6dbf51bf808fd3f0187095af43f0149f788;
mem[99] = 144'h06a7f0daff4ff2ebf783009b0b96f42f02f5;
mem[100] = 144'h052aff200389f58c04ba0da2018108900161;
mem[101] = 144'h013f067bf3bdf1f3f41800a0f25109cafdbf;
mem[102] = 144'hf5cdf8e9091608b40601084eff9ef61cf37e;
mem[103] = 144'h03c30d43f4450f1af62a02a0f05bf7f1fa2c;
mem[104] = 144'hfb0efa51f3aa0dd9fca00ee9fccefd400e77;
mem[105] = 144'hfda70c81f60a0a9e04fbf2ba0f9a034cfd53;
mem[106] = 144'hfc54fdc103a90032f99afa3606d7f2d50d2e;
mem[107] = 144'hfe82f153024bff3af96e0a8cf53e0fdf06b4;
mem[108] = 144'h0ac2041c00bb085b074f092b0eacf779f0cd;
mem[109] = 144'hf63ef0c902f6f2c90523fe0cfb75037b03b5;
mem[110] = 144'h05680cf30036fdec046909e10608f4e40550;
mem[111] = 144'hfc45f7290e8efdc7fb0c0e4502f4fc5a0f96;
mem[112] = 144'hf9e80ecffd40f1cef097f4bb0df90b98f3a7;
mem[113] = 144'h0eedfbd2f64dfdd505680a54f5b4f8a5f008;
mem[114] = 144'h07bb078cf44e0015f69ffffe0cbdf1a4f4df;
mem[115] = 144'hf66e08cd015909b5f13b0192013bfc50fdc7;
mem[116] = 144'h00190a30fbfffad7fdeff6a908d7fa65f5a3;
mem[117] = 144'h02220eb4f56507f0008ff85f06ed04d9f6fc;
mem[118] = 144'h0fb205ecf800041400c20a170f43fbf309c5;
mem[119] = 144'hf732f0d5089309d1f6300dce0572f1980806;
mem[120] = 144'h06a9ff9afb280719067d0b430e96f3570ecc;
mem[121] = 144'hf52909fe0977f3af09200db3f6dffef5f822;
mem[122] = 144'hfc38fb91f9070261f12809a4f5580e580802;
mem[123] = 144'h0258049a0d06f5a80852f865f626f9f0feeb;
mem[124] = 144'hfe6f0b56f749f7f603e6093efa26ffe8042f;
mem[125] = 144'h08880248001bf84100690083f13b0b50f976;
mem[126] = 144'hffdd0054fac1fcc301fbf32cfb58f2f4f5cf;
mem[127] = 144'h0bd9f09bf9e507f0022f0eeb0baa06b6f45f;
mem[128] = 144'hf8b9f7e8fd47f1ef031cf229f02000cd020d;
mem[129] = 144'hf41606f10d0ff04cf7b30c9ff317fa08f870;
mem[130] = 144'h078f0646f095fd25f11d0070f109035afc5e;
mem[131] = 144'h0f7bf64a0b5e0567f0480663f9ecf02504a4;
mem[132] = 144'h0c4509e904900fb2028bf464f8cb001e02bf;
mem[133] = 144'h0b9907d0f5dd0037fc9b0acff831ffe60530;
mem[134] = 144'hfdd5fbe6f2a9f505fc24f9a40c57fa8002d5;
mem[135] = 144'hfdc306100f2bf37e029c0be600d1fb630c25;
mem[136] = 144'hf138089c0b1ff7f9f3b50501f2eb062a0435;
mem[137] = 144'h0203f2c7f441025dfda2f0fdfb0ffdad0ff3;
mem[138] = 144'hfaa4f87407f3fd7609bdf996f0270ba60fc4;
mem[139] = 144'hfad3f7da0f37fd8ef500022cfe66030cfd44;
mem[140] = 144'hf882fe0fff92f55205dcf3a10e80fb16f91f;
mem[141] = 144'h04e9f477fcd6f4a2f1ef07a50767073ff371;
mem[142] = 144'h0076fe430695f203f544f4ff01ee02ff09f1;
mem[143] = 144'hfa780edefaa8fc4efd69f143fc5df65ff9fe;
mem[144] = 144'h06def321f616fef2fc52f2b6f2f60e6104fe;
mem[145] = 144'hf90e08f30653014307fa0e1bfb4afb9b0e86;
mem[146] = 144'h0edeff480844022df91d037e0114f53bf334;
mem[147] = 144'hf1c80c99fb7206e8fcf2fcaf0e7fefee00ae;
mem[148] = 144'hf13805df0a17ffe002b60215ffc2f68204af;
mem[149] = 144'h05cdf3eefbd30b39fa24f99500980f19f281;
mem[150] = 144'hfb31f2980434f2c504a5f8d7fb9f067ff7be;
mem[151] = 144'h05510eaaf95cff050900ff680f13f40bfdd1;
mem[152] = 144'hf8b6f662fc78f81402d0f4e2fcf70acefc9d;
mem[153] = 144'h09130dc60a79f746f2370a4bf6b1f5ee0341;
mem[154] = 144'hf163f0520c31f590fe4ef4e40af801bd09a8;
mem[155] = 144'h09600bdb08f6f6eefcf1fb12fe6b00900395;
mem[156] = 144'hfab9f1fbfb33fd1d09c4f770f7f30d520021;
mem[157] = 144'hfd7c03960642f8fffa600116f9a60e3e0792;
mem[158] = 144'hf1780283061700e9f3810435091401510860;
mem[159] = 144'hf409f54f030df622fabf0360fa2608330c18;
mem[160] = 144'h07d8017202b30061f6a5f60801b4fe8ff78a;
mem[161] = 144'hfc3d076e00020a7704b2078c046f040f05b3;
mem[162] = 144'h012f0764fc17047cfe8b089d09390ae0006a;
mem[163] = 144'h0d78f8d9fc47fc970d1df93701f20619015c;
mem[164] = 144'hf9d5fb80f5bbf7960d28f7fdf530efbdfd8a;
mem[165] = 144'h061ef0230d280abd04d8009cf589f22e09fd;
mem[166] = 144'h0d9c056406cdfbeef4f6fd0b0b240c1404ee;
mem[167] = 144'h0146f6ff0028fc01057ef47c0b32f334068a;
mem[168] = 144'hf96b0d4d02800de5fc56ff8ef454fc84faab;
mem[169] = 144'hf0ac0532efe5f179f656fa86fabcf410042c;
mem[170] = 144'hf65c00e9057bffbb061ff5a20033037ef17e;
mem[171] = 144'hf669fc7bfa250881fb5bfb9c07e1fbbb05ef;
mem[172] = 144'hf88cfd730bc5f63407ee0e6300110c61f6de;
mem[173] = 144'hfc740130eeddf6f503b3f0a90c65fd0d025f;
mem[174] = 144'hff67f9b9ff24f482062df83806b507bef0f2;
mem[175] = 144'h092ff6650183fd4af164f3b60f050a72f95b;
mem[176] = 144'h063508010dd50623f2eff73a0da0f20a0d5c;
mem[177] = 144'h0f98f1c606a2fb510687f287f06605feef6f;
mem[178] = 144'h0e9d09e5f7510bdf0f86f93ff93cf635025d;
mem[179] = 144'hf339fe9400a104a802680ef00ed800f3f360;
mem[180] = 144'h0aebf5410515f2910857fea104b5fd3e0901;
mem[181] = 144'h0cce0366f265f35af585f6970f730673f51e;
mem[182] = 144'hff8af1e5f2ebefae0e64f26008f0f77f0252;
mem[183] = 144'h09d2092e047007aaf79909d10f6009e9f34f;
mem[184] = 144'hfcb70ed4f4a8f236fff0010a0ea5f799092d;
mem[185] = 144'hfdeb09f707e2f7dd05d6fbef0c4a06e404b0;
mem[186] = 144'hfd1ef5c10924f7050b180c6e0a23fced0ccd;
mem[187] = 144'h0f7a080e0739f9e70758faab0cd9f155fe5c;
mem[188] = 144'hff19fbef02b50e54fe890a7afce80b24fcd2;
mem[189] = 144'hf7b8ef8afe2804970751ff18efd6f27cf4b0;
mem[190] = 144'hff09fea10ccdffdf0317fe980b4ff93ffbf5;
mem[191] = 144'h0448fa52fb0e0c64f06e0f96ff28016cfdef;
mem[192] = 144'h0f41fa7801fe0baf011105730475054402d9;
mem[193] = 144'hf615f3ba0c9bfb2b01ed011b07df0e17fe61;
mem[194] = 144'hfc060439fa67ff72f3b4f04a082f074afa9f;
mem[195] = 144'h0aef0868fda9fef1f1cffaa0f1d6fd8ef1e9;
mem[196] = 144'h0d150a7efb76f3e90ed009b7f1abf9e2035c;
mem[197] = 144'h0bd606470ba60be1fa8809730daaf42e0e52;
mem[198] = 144'h01f9047c07870643f820ff34fb680f83f88e;
mem[199] = 144'hff2a0f55f6c00b600a35f5990eb2f90d0c89;
mem[200] = 144'h0d270156f655f9befc08f14d0036ff2b0bb6;
mem[201] = 144'hf193f6f2f54bf92b0868f138feee064af440;
mem[202] = 144'hf94e00320d5000f4fa87fbe60995f506fccd;
mem[203] = 144'hf1f60326f4bc0ebb0d570d2b0c6c083803b4;
mem[204] = 144'hfc4a0f970f600430f0280902071900e3f5e7;
mem[205] = 144'hfbf604caf9fe0014003efedb02f20696f7d9;
mem[206] = 144'h033201c5feec0f530e9ff36403ce03b60199;
mem[207] = 144'hfecbfccdf53cf3e0ffebfab20009f9920f55;
mem[208] = 144'h0cfff9770cf80a09f80bf333f9d702a509b4;
mem[209] = 144'h02d90a83f6aafa7ffad803030d8e0191f5cf;
mem[210] = 144'hf63df82f0de3f9c4fc36f2c0f00df2560400;
mem[211] = 144'hf8eaf298ff750928052cfc080d9d00790cd3;
mem[212] = 144'hfd5c0f090b41f0e1f7730d00fb0d0d20f53b;
mem[213] = 144'hff7af30df2e30ae70b8809fc02d8f3110d89;
mem[214] = 144'hfa6f09610e4d048cffdcf7720f0e0134fa24;
mem[215] = 144'h0335f21ffa140caf014cfb070491f3aa0169;
mem[216] = 144'h01b70219f227fd54f859fa5d00fd07850808;
mem[217] = 144'hf579f6890d1106baf388030bf23c0bc40478;
mem[218] = 144'hf724fffefbeeef91fd58002ef97cf847f197;
mem[219] = 144'h04bb04b002f009cbfa47f03ef2d0f44fff83;
mem[220] = 144'hf2560696027ffadd0c08f4e20d59057ff18a;
mem[221] = 144'hff20f34af8b403ee005df506079af8410984;
mem[222] = 144'h0a22f9d0f4b9048af872082a08fef3280d43;
mem[223] = 144'hf847f325fe73fdfe034404a20256fc660ad8;
mem[224] = 144'h07cd02580e78fb31083e0dcd095e042af2e9;
mem[225] = 144'h02f104aef159ff13f027026df4140600f1f4;
mem[226] = 144'hf3f1f18af645f678031efa3901990dbcf9f4;
mem[227] = 144'h045defd4fd250360f20f0394fc9bf78f0735;
mem[228] = 144'h084cfa70fd07f0930a48fe7609e10dc30a91;
mem[229] = 144'hf8160ec9f492fd9007d901f307fe0779ef62;
mem[230] = 144'h0dadfdd101d7043106a0f66ffa70fa27f831;
mem[231] = 144'hf7910b68fb3af475fb360142f78c09bcf2b4;
mem[232] = 144'h0726fb75f6b9fb70f01602930c5e0538ffb1;
mem[233] = 144'hef110bdc0a8204590002f185f73af457f1f0;
mem[234] = 144'hfc3a0859f54df878f2d3fbf5fc6af132f195;
mem[235] = 144'hff7c0ae0f6c30ce4f2c8fd1d0e350d030bce;
mem[236] = 144'h0e82081203bdf888030aef97080e093f0238;
mem[237] = 144'hfec0febb0edd03830d38083af01b0051f0de;
mem[238] = 144'h0db70dca0e860299f0c5064ffb68ffff0832;
mem[239] = 144'hf9ae05fcf0960210fe8e025201bd0b3b0f37;
mem[240] = 144'h00a7ff2df8a907b4fcc909bd0cacf0bef509;
mem[241] = 144'hf24ef8ca094b01ecf0f40c08084f0a4cf584;
mem[242] = 144'h0a52f9c80146020706620215f90c0f20f361;
mem[243] = 144'hf8fd0215f83dfb29f76efefc0c9e0ce1fc45;
mem[244] = 144'h05cf0b2df27303370a67f8c1f0f6fbccfb43;
mem[245] = 144'hff02f88a04effa98f1680f98017007d00b95;
mem[246] = 144'h0d21fbb7f4eafe0ff3380b570a6a00290b36;
mem[247] = 144'hff820479f203f934f6e5f84607dbf3150bda;
mem[248] = 144'h0a200daaf7e7f84afbcff93f07c804f3fa55;
mem[249] = 144'h0d49fb78043402fff52c0c2d0126f11efb66;
mem[250] = 144'h0b23f97bf40afe0d0978fabf09920b1403af;
mem[251] = 144'hf3080f8af331fc94ff020d9e01b6097f039b;
mem[252] = 144'h0a3bff6e0d95056beffbf8a30c54f086f6bc;
mem[253] = 144'h0344fd590f88fab7f3a3f3adf770fa47f59b;
mem[254] = 144'hf2e1035d0f83f7ab0a6308ce0fa40a2af16d;
mem[255] = 144'hf626fb380a19f4dbfec6f3780637f2c2feae;
mem[256] = 144'hf3a7f7d7073607090ce40a1202b602cdf5dd;
mem[257] = 144'h0640f679f100f4390a8707adf62c0a2f088d;
mem[258] = 144'h064d0faa0ad6fa1afcbf056efbf104fff099;
mem[259] = 144'hf9a3f145096afd87f048f3cf094f064bf80d;
mem[260] = 144'hfd280752f39df57306f6067c04cf03890ae5;
mem[261] = 144'h075ffce70690f93bf8860c9b0acaf694fbb5;
mem[262] = 144'h01150950fbb20ac3f3da0e75000def600df5;
mem[263] = 144'h05ac0ecbf3bcfe160a9ff108f4f60408f16a;
mem[264] = 144'h0c9707da0d1e062f0eaa0a860a49ffa2fa27;
mem[265] = 144'h0becf6fe06290accf70df046fe1a0ea30bf2;
mem[266] = 144'h0409f83004030a170544ff1907b7f976f315;
mem[267] = 144'hf43e01fb0a61fe70f02701d0fc9aff51fcee;
mem[268] = 144'hf08ff57b08c90b920b89f42e06110f0bfe22;
mem[269] = 144'hff5ef72ffd040aa8f8b7066d01850e1cf07a;
mem[270] = 144'h0955f0b703e0f335018e0e0efe5cf9920175;
mem[271] = 144'h08aa0849fc57f4d0fb21070cff44f3a407b3;
mem[272] = 144'h05b00613f185f103fef1fb9df601fbf50cfc;
mem[273] = 144'hf5990851f23c0fac0674f486035df5780e84;
mem[274] = 144'hff37f9b9f89dff16fb77f3bffbb60a37efe9;
mem[275] = 144'h0157f47af544f7b3f3c8fb29f978fb4507db;
mem[276] = 144'hf3d1fdde056bfbbdeff30c2005f1f58ffcf8;
mem[277] = 144'hf1f2efaef83b08d70d13f506f777f8a0f2e0;
mem[278] = 144'hf8d80716060ef7690a49fc3f0711f4ae0269;
mem[279] = 144'hfa8902da038402c3f8f1f9d1093400040c66;
mem[280] = 144'h0e5a06bffa2d0e4404e7fb3cf55a00d4f6c0;
mem[281] = 144'hf421ffda051b0b1a05390616f6fff5820e36;
mem[282] = 144'hfc840375ff59fcdc0ceb07970cbc0231f835;
mem[283] = 144'h0770056a07e9f02ef5490a490d980f6af4bc;
mem[284] = 144'hfd290beaf2fdfac5f976feffefbf044efeea;
mem[285] = 144'h0e35f7c408280187028402cb0bb107b8fb9b;
mem[286] = 144'h0b1bfaa5f844f7460d3b08760dd3f7e9fe76;
mem[287] = 144'hf8eff8d5066ff2b607db09e8f547fbd3ff6e;
mem[288] = 144'hfdc60f0100d101e1f69605c206cb08df0b9d;
mem[289] = 144'h0969f38bfe79f9a7fe49f14efa8af4b8f1f4;
mem[290] = 144'hf8c3f0ddf9c502340d74f2c9f9e10e93fe8a;
mem[291] = 144'hf4ae0510f948f87ef615fa8b0f0cf3c10021;
mem[292] = 144'hfd910c1ef7370836fb1e069b0a630a78f6d1;
mem[293] = 144'h0cd1f8f60c9c0e93f1b2fd34f2b3f4aeef0a;
mem[294] = 144'hfbf609250d5203bff52d08f2f47ef350f79a;
mem[295] = 144'h02f9feaff1390b0002fbf7470145fcb800c2;
mem[296] = 144'hf489f5b7f3260b9e0a76f20bf5b701acf172;
mem[297] = 144'hf856f88a0ea209e10b7b0701007104b502f5;
mem[298] = 144'h01140b8d03720651f762fd70014ef6d6fc75;
mem[299] = 144'hf2a1035f05dff750f9dbfe660a96fdb3f5a7;
mem[300] = 144'hf4250b770bd007cbffbd0b21f8dbf7f90e3c;
mem[301] = 144'h0db90763f40bf28d01b8fe850d67f5770a92;
mem[302] = 144'h084e053b08910ac000aff45e0633024b0210;
mem[303] = 144'hfebdf8190389ff46f82505f402a9f5fb03a6;
mem[304] = 144'h0833093ef834fa6bf304f29502e0f6c00a8d;
mem[305] = 144'h08470087feaafb31fc1707b3041f0d49f55a;
mem[306] = 144'h0b1509eb0085f2930bfcfee1faebf7890b92;
mem[307] = 144'h0efff7bd0abffa38fd70f452fd15f4e90d32;
mem[308] = 144'h0ba9f1dff429fd110b42f99afc1ffb7504e7;
mem[309] = 144'hfe8f0f0f0f4c0baef680f8d7f2e7f240fa2f;
mem[310] = 144'h0468069c08f6fef1074df601016f090c0b20;
mem[311] = 144'hf8f409640599f22f06c407210958f8ea02de;
mem[312] = 144'hfc290f3bfe380675ef9a00ac0c5f04fa0b28;
mem[313] = 144'h086afce3f0e5ff82fcf6f8b3f04f0e740d07;
mem[314] = 144'hfdb4f470f76df07cfc95ff850dde0747ff93;
mem[315] = 144'h0b2efe55fab6ff47f2b2f0fe02970d1bfe20;
mem[316] = 144'hf5650640f7e4f809f2bff5ef02a100860cbf;
mem[317] = 144'hf4840cf10695079b0c1d06f2f2ebf87e05bf;
mem[318] = 144'hf829f60ef71ffac8f909036309a80accfc52;
mem[319] = 144'h0e9305adfaed0f3c0e1606a50327fb52f8bd;
mem[320] = 144'h0f28f31307e9f0330c380e37f72a02af02cc;
mem[321] = 144'h0065f57f000ceff0ff4301dffd77fb610e68;
mem[322] = 144'h037f0e92033df6c107a0f077f43e0787f23c;
mem[323] = 144'hf6bb0a070f8f0c83f2d80403f856fcbe0385;
mem[324] = 144'hfdf1f7720d15074efad20b4afcce0bb2f600;
mem[325] = 144'h0291f7a1ff04ffcf0e76054df67df1fc0302;
mem[326] = 144'hf041f086065dfa090054ef760d10f58507cb;
mem[327] = 144'h04f106d8080dfe3f044800e8037f04130aeb;
mem[328] = 144'hf11f0350061b0c1b0f9af34f05720e450deb;
mem[329] = 144'hf443f40cfae6fb4e05c0f29205700927f468;
mem[330] = 144'hf80ef1d20f4df204f4300450fff4067001a9;
mem[331] = 144'hf2d9ffe7f4f9fd530cd1f7420e91f337f1ed;
mem[332] = 144'h0af5f00e002202780171feeb0c64ff72fd78;
mem[333] = 144'h0667f151fa72f62402ca0cb4049a0d080c31;
mem[334] = 144'h0863000b07d5f3d5f55101a70cad042a078e;
mem[335] = 144'h0d20030904d90b5700eb0fad09f3011a0488;
mem[336] = 144'hf3640c430de8f08ef6ef039a020a0ac40b2a;
mem[337] = 144'hf430f080ffad0f46f3460d5e0188f8a60797;
mem[338] = 144'h0789fba7fcaff1e009ae0151fdb1f4b80681;
mem[339] = 144'hf220f411f9fa08c3efa207c0f033f2d40783;
mem[340] = 144'h0ab2ff5e0006fe1703d9fcf900c7efde0837;
mem[341] = 144'hfbd207090127fddef5710e11f215fd29f369;
mem[342] = 144'h04120326062bf199fcc6f6b00c70f550f6c2;
mem[343] = 144'hfbd1f8f5ff690dda0a830a320ac90e80f20d;
mem[344] = 144'h04d701e5f969f8b7f01ffd67f2690134f0c6;
mem[345] = 144'hfe22fbac0c76f530fc2f0e02096c075aef14;
mem[346] = 144'h02cf0b34f0ff0cfe0cb9f99b0382054a08b2;
mem[347] = 144'h0cd905bb0ebe0f9e08ec0608023ff45ff903;
mem[348] = 144'hffacfe6ff06af8e304dbf8eaf5b8fb7606b3;
mem[349] = 144'hf4570e8bf226f7c2faf80da3f04507bf065c;
mem[350] = 144'h04c2f425fbc607fd0d920849f6fcf17a0d3d;
mem[351] = 144'hfa2cf5e9f57bf332f742f8d9fca60e88fd94;
mem[352] = 144'hf86e0dccfb08ff060e4ff827f253f5fff9fb;
mem[353] = 144'hfb4008a10839fb7af5bbf9f1042affdafd3f;
mem[354] = 144'h088502cffa4a0781fff8fb2a00b6fd54fce2;
mem[355] = 144'hf1c0f5d7fea4f21e0dc7060ff376f708f18c;
mem[356] = 144'h06eef89ff65004f3fb3e0f91fa02f154fb63;
mem[357] = 144'hfd220da3f493078bf2f709e2fbc50708fa64;
mem[358] = 144'h076d0b4d0ca2f123068bf4b40c34febb0972;
mem[359] = 144'h08b2026b02fc0c020b9803960855f62af1cf;
mem[360] = 144'hf43b040807d70e63f879f7ab0c3af4040835;
mem[361] = 144'hf5dd095af1d8ff8d0a9c0aabef43faa5fa45;
mem[362] = 144'h03fdef6dfb58f0fe09f5085801fef48b0773;
mem[363] = 144'h06e30d63f41df6d8fd81023f0d59fea5f569;
mem[364] = 144'h0535fd5e088802ab01d5077ef9c506a3fae7;
mem[365] = 144'h01fd067ff54f0ef4078cf557f4d2035cf439;
mem[366] = 144'hf56cef98f617fb960200fa8400bcfd8b0a26;
mem[367] = 144'h02b1fe7b0ce3fc020574027cf232feedfd16;
mem[368] = 144'h000c069302f2f73c025a0bfef774099703f5;
mem[369] = 144'h0299f1e207cc0888017f0af9092a0b0affcd;
mem[370] = 144'h067efa75f9ecfe3df6050fe2037cffc0f568;
mem[371] = 144'h0e8ff6650c51ffa6f7170c89081700a6f135;
mem[372] = 144'hf82cf33ef8c900500bbe0f9afaac0027f520;
mem[373] = 144'hf1e2f9ea0fc6082f08ccf37ffc9bfb4af039;
mem[374] = 144'hfad70e110184ff3e0a45f6eb0781f059f0d9;
mem[375] = 144'hf4140f06f10408670d9e0efbf01afdd8ff43;
mem[376] = 144'h0dd3f2a3f01ffb37faef053b01da0227fd23;
mem[377] = 144'h00350e780524fd0afb010c75f95100170f9d;
mem[378] = 144'h0993023f06ba04130875f618f6600703036e;
mem[379] = 144'hf2f60ecdfb8dfa8af87d0fb8fb11f081096c;
mem[380] = 144'h0c3cfbe2fa86078c00bb0f87f3aef3a6efbb;
mem[381] = 144'h0954fa2001abf9abf41f0640ffc20715fd9f;
mem[382] = 144'hfaa9061c06980025f11806360e63f1530dd4;
mem[383] = 144'hf4b5f5cef9f5fa3af76007f3f51ff0f6f2a3;
mem[384] = 144'hf8d30a4005f4041bf253f6c7fa21029af9ec;
mem[385] = 144'hfeb2f3d0fde90f6f0171f9d9f2daf71507ee;
mem[386] = 144'h058e0607ff32f53defe5f58e071a007cf0b8;
mem[387] = 144'hfd5ffb13004b039b0424fd600dd0fd520967;
mem[388] = 144'h044c01de0828045af3c9fc63013a0b030876;
mem[389] = 144'hf2cff65efab0f406f0250067043b0503094b;
mem[390] = 144'hfca8084105f2fe29f7240f00fd3afba8ff0b;
mem[391] = 144'h06950654f986f761f786fbba0d83fc7b01c8;
mem[392] = 144'h0a2808cbfed4fe29ffa405c70864f2c701c4;
mem[393] = 144'hf29d0e44fce309faf868f63d009ff5faf7bd;
mem[394] = 144'h08890cbdfda5fabfff320dbd0b2af333fce8;
mem[395] = 144'h0f50f0710f07f1450f2505bffd180e0608e0;
mem[396] = 144'h00c7fb770145024901fffbf30900f7e4f56a;
mem[397] = 144'hf7b2fc95063bfbfafc040289057c0406f1f4;
mem[398] = 144'h0ad1016f0a09001dfbf0f66bf120f7edf246;
mem[399] = 144'h0d2900cc02db00fff3ea018afc22f68c0467;
mem[400] = 144'h022408c1fab10142fabbf53ff53c07f3f8fb;
mem[401] = 144'hfddf0a740f4904cf032403f80998f745f3b7;
mem[402] = 144'h0cde02830b7ffa0df07c03940877028df4ec;
mem[403] = 144'hf7910ab9fa14f2b0f19cfaa9fd8ff31dfa0d;
mem[404] = 144'hf05005a9f06201ed0ab1fe0602fbf8c8faad;
mem[405] = 144'hff2af6d40603059101ebf5fbf35ff5be00f0;
mem[406] = 144'hf262086d07ddf491fa46ff0e07490d69fd53;
mem[407] = 144'hf201042afc07faf80231f183f6b5fd400f32;
mem[408] = 144'h06d90f1bfaee0dfa054df3110912f5ccf63e;
mem[409] = 144'h0f51fb62093b004af2200c36018afc0b03cf;
mem[410] = 144'hfdeef5f604160c6b0e9301e9f4b40ce40fe5;
mem[411] = 144'h02faff79f881ffebf7bef4a709b0f0ae0384;
mem[412] = 144'h02270242fe11f5a9fabafc52046003d90dd7;
mem[413] = 144'hf533fdc304bef59207640be3f7150792f736;
mem[414] = 144'hfff400d002caf4edf90b0454f3db0e7af295;
mem[415] = 144'hf83efaf7fc280420fb48f792f70ff5b6fef1;
mem[416] = 144'hf7c1063ffeb0fe3009edfccdfc8b08edf200;
mem[417] = 144'h09830c330677f8d2f2a2f41801e50b680bbd;
mem[418] = 144'h0e2c0f25f5230dc5f659facbf0b6f819f901;
mem[419] = 144'h096405e3f26703e70704f8bafa36f9fbfcfa;
mem[420] = 144'h0f5af81ef5b5f46708ba017cf852011e0233;
mem[421] = 144'h037e079cfa040097fd6908e1fd0402c60e9d;
mem[422] = 144'h0b840f40075af5a2fe39030bf5d30af908f8;
mem[423] = 144'h0829f0a8010df482f3a502cb0243f1c00c2f;
mem[424] = 144'h02e3f800f7c9098505d802b9f1bcf1910bd4;
mem[425] = 144'hfa63ffdc0ece0c100336058dfda2f6ebfb88;
mem[426] = 144'h0163049803df0caff62ffbf7f92b010e06da;
mem[427] = 144'h0c910dadf9130947f91ef7b40129f51e09b1;
mem[428] = 144'h040cfb0106c907bdf139f0bff110f7cbf166;
mem[429] = 144'hf278f6e001c1016e04b3f0560dccf420f0ca;
mem[430] = 144'hfd8af0cafa490d7cfeb5f3cdff610138020c;
mem[431] = 144'h09390e5a0bd8fe79ffd608f0f17afeadff70;
mem[432] = 144'hfaef0e6e0e7501d605800b250392fc75f327;
mem[433] = 144'hfc660117f8d6fc74fc2b0f69fec2f03f047c;
mem[434] = 144'hf3bb09f5f317f4330117f353fc250e8efcb0;
mem[435] = 144'hf51cf093ffa9fa2a0cfaefda0572f274f173;
mem[436] = 144'h06b5fe79fdadf9ebfbee0e6f0f9ef6d5ff3e;
mem[437] = 144'h0d19f3feff09ff9e0b750dd9f8f8f2df08e8;
mem[438] = 144'h0ce206610ac20a1500a4f329f8e103a0ef2b;
mem[439] = 144'h06e60e500780f67c016f0245f984019ffa6d;
mem[440] = 144'hf1c2005a03c5049ffcb3f6ecfeaf01980365;
mem[441] = 144'h00c8074b03a1fa1603ddfeb7f0aef6f3fe74;
mem[442] = 144'h0899f2370cd7035df061024f0564f711052e;
mem[443] = 144'hf847fd22024efce4fe21f334ffdffff1f347;
mem[444] = 144'hfe88f7c7f4dd00f1f3d5f05d082f06f4efc4;
mem[445] = 144'heff9f23b09bffe6b032d05eff93f0981f475;
mem[446] = 144'hef71fed0f580fbe10a38ef10fb30f4560bf5;
mem[447] = 144'h0a240a93f521f4d804850d1b0051fe45fcbd;
mem[448] = 144'h0592030af50f06650e73fef8f4b2f6fc0580;
mem[449] = 144'h03710487fa42eed2fb7f031a0fee00b3ffa5;
mem[450] = 144'h0f90f7caf6240f2303d9ffb9f782f77c07ca;
mem[451] = 144'hf3f302d50a5900640b6708ce0e160a38f11b;
mem[452] = 144'h06dd0c5d0e3af1f80904f8230c3c0d13fec1;
mem[453] = 144'h05b00b57fb7c037206770b58fa22f3e6044c;
mem[454] = 144'h05e7f0f6057bf6b202b9f4c40190f03a0344;
mem[455] = 144'hf70cfc390f490c20fb63fc870feaf93cf15d;
mem[456] = 144'h09ddf9490e0ef6d90793f33304d9f01df2e9;
mem[457] = 144'h0f97fc03f3d1fc5d03a0002bfab40ab20c0e;
mem[458] = 144'h075d0bcdf3540dbbf470fd98f780f70cf55c;
mem[459] = 144'h0630f829f81ef3c3ff9efd68fe5bf35d0a28;
mem[460] = 144'h0757f9aef08a0f28ff90f75d028ef7ebfb47;
mem[461] = 144'hf558f5540ea3f79efa24f284085ffa030418;
mem[462] = 144'hf399fdd60830fece085a045806edf79df359;
mem[463] = 144'h0b5dff090514f8a908bafe910f2505350317;
mem[464] = 144'h04b905780cfd01ccffdd0ec50e510552fcaa;
mem[465] = 144'h0389fa980c19f65f0e7609690531f2e4f173;
mem[466] = 144'h0235fba10074ffbbff5208effd61fce8f2e3;
mem[467] = 144'hf4450734069df41ff566088c0d4af7ec093d;
mem[468] = 144'hfc38f3640996099f0e7b0f2a0dc8f44eff4b;
mem[469] = 144'h080c0b82010ffd89f4eef49ef137002cf9cd;
mem[470] = 144'h09310aacfef90732f781f0a7f2cd0e3301ef;
mem[471] = 144'h06870e64001b0d94fc68f323fd84f19efd50;
mem[472] = 144'hfd3c03cbfdc6f63bfe5ff4e005a7f2f9fa3e;
mem[473] = 144'h057301f8fbc3063cf23affa4f225f24af665;
mem[474] = 144'h0452fa510bbd0dedfacf071b08d2081f0019;
mem[475] = 144'h01880816f325fd57f89b03ebfcfc03ed050e;
mem[476] = 144'h07bf0aa4fc7300eb055df616ff970500ff64;
mem[477] = 144'hf69002000aa4f71df2cc0822fe900ac10b33;
mem[478] = 144'h081ff0b1f8a2f1a3f6480ce8fd9df575f1c3;
mem[479] = 144'hf167f4a8fd1606c60fc4f1610c75f5b3feb9;
mem[480] = 144'hfd640e940fa7fe50f21df6f1f11bf3580510;
mem[481] = 144'hf5c9face0d60f9a400bdf5ccf8500b82ff3e;
mem[482] = 144'hffaa0c65073302a1fcb709edfd1cf511099b;
mem[483] = 144'h02a5f4de0ca9054602adf156ffee02b8f794;
mem[484] = 144'hf4a8ff0f096c08abfb81fdc0f3250f1defd0;
mem[485] = 144'h05a4f798f8a7f574f1ec0760f01bff4b06dd;
mem[486] = 144'h0dbe0c660e9f0402051e0b4e024ff49c07ba;
mem[487] = 144'hf983fb670693fa18ff26f71700cf07f506fc;
mem[488] = 144'h07f5fe72054af875fd50f67df2b20beef927;
mem[489] = 144'h08170b29f09000c8f4d30584031df7c50a19;
mem[490] = 144'hf6a3fe6a071b014608f4fe91f967f980ff18;
mem[491] = 144'h0707f5d3097d092bf41f076106d800680178;
mem[492] = 144'h0b8affcdf3f207d40707fb2d00fb0a79f4c5;
mem[493] = 144'h0f4ff38ff4f60a7df5f1f844090cfab50344;
mem[494] = 144'h02d201c604e9f471046106b80346fa60f428;
mem[495] = 144'h064b0136f6c7f4acf64c0ae8f417f485061e;
mem[496] = 144'hfa3e0aef0343f063ff66f7f708ba01b704a6;
mem[497] = 144'hfa52fcf7f416f3a8f7a4f321054cf801f54a;
mem[498] = 144'hfa60f8490da5fa7003dd0f8208f1061002d2;
mem[499] = 144'hf764fff0f0ff049a00baf57ff94409b40196;
mem[500] = 144'hfbdcf3a5038ff1f6eff3f3410c47fa4ff917;
mem[501] = 144'hfd8d07a2f441f6db04c0f91e0417fb5c0978;
mem[502] = 144'h0278fd40fc1c097c0d490b1dfa1df6c8029e;
mem[503] = 144'hf7cbfbb403ebf04608b0f8fa0f49014c0dc4;
mem[504] = 144'h0fab058303e1ff19fb690cc308c6f21504b7;
mem[505] = 144'hf442f8130bcafbb70da604b3f053fbf50f3d;
mem[506] = 144'h077cfe9f0af20b60f24c08c7fdf90c07f8de;
mem[507] = 144'h08070309f3540ef40f9c09c70d900ec8fdf6;
mem[508] = 144'h0cf5097af5530c97fa5bf4080490f26d0a1d;
mem[509] = 144'hf64b03a3f4a0f6bf0e190ee2fd15020d048d;
mem[510] = 144'h09fafcf1ee2e0763f366fe4c0151f72f04f6;
mem[511] = 144'h083fffeff37df3e1085bf55bf215f456f1a8;
mem[512] = 144'hf75b017bf143f6ee090804050d4908990582;
mem[513] = 144'hf5320ebd092bff1df81bf801f9350981f402;
mem[514] = 144'hf488f3abfcd00008f02707f1fb8f0391f817;
mem[515] = 144'h0a8fff6e05b2f339f4f8fe750c6903fff704;
mem[516] = 144'h0dbd0c5502e3f481f7ddf9a505660c680816;
mem[517] = 144'hf18af7ac0751051b0b64f17ff17f0a98f149;
mem[518] = 144'h0615f13f0a8df593fd50fb10f0db0689fa58;
mem[519] = 144'h0e79f168020efc4dfc3a0541fdb108dd0bff;
mem[520] = 144'h015f00bcf6740bddfdf9f49ff0db0d70f519;
mem[521] = 144'h00ebfb0df0b40f3f00350188fdb1fdf2f63f;
mem[522] = 144'hf092f5270c61f79cf055fab70dc5f32f0eb7;
mem[523] = 144'h0c2d03a2f9d0f89805f0038cfdb2f8dcf887;
mem[524] = 144'h042bfbb10b4407a8f5ef04fafa57f09efe85;
mem[525] = 144'hf64f04030961fa630136f77efab80304fddb;
mem[526] = 144'h0ee1f1a2f7ea0d5902ac00b1fb5af611fb9d;
mem[527] = 144'hfdc2fc5c0e0e00f0f52002b60156fb0a05ac;
mem[528] = 144'hf798fcf0fbd5fcc6fec10b43f0b9f567020b;
mem[529] = 144'h00c7f0f30ad4fd1af273fd88ff4bfe20f2ea;
mem[530] = 144'h0fd7fd5d06a5f34606c7fa2df42c0d88075a;
mem[531] = 144'hf05df0fb091205a503d405e009ec02c20cec;
mem[532] = 144'h0bbdf1f20048f284fcdb0ed3fa14f0bcf7db;
mem[533] = 144'h0c5cf01ff324f8290a43fbdcff8c088af611;
mem[534] = 144'h0a62fca7fc72fad7096102c5f687f797f562;
mem[535] = 144'hf90a0b79f309fd26072f0275ff82ff980fa1;
mem[536] = 144'hf285f9810d460f680e1ff25afc69f6c2fe60;
mem[537] = 144'hf9a9fae6010d06eff68401bef3faffbffcae;
mem[538] = 144'h0d74f41ff875fbd60d89faddff77f41efbfa;
mem[539] = 144'hfa9eff0bf5e90850f2960242029a0843fae3;
mem[540] = 144'hfe0df26afbbb0dfdf9a90c8f04c2f14af904;
mem[541] = 144'h08b7030afd030801f70cfdbcf37e07dbfda7;
mem[542] = 144'h0a21fe290e22ef7d040e0345f76604080167;
mem[543] = 144'h0697f05c0f62f31fffa4f232fc70f109050a;
mem[544] = 144'hfd4100530965ffcafe170adaf8ff070ef17a;
mem[545] = 144'h0822fa9bf79e056d09b705720528f6f9f32f;
mem[546] = 144'hf17ef5f6f7edff42fdd704d6045b00ef0a50;
mem[547] = 144'h05eb0153f5810be80aa7effaf6e704e1f9dc;
mem[548] = 144'h08ea04900769fb7ff092f5010e1d06e30bd9;
mem[549] = 144'hf472f07cf12d0c2ff8640cdff588f5f6f75f;
mem[550] = 144'hf9f608f1fb9f09040519048208b50d5cf524;
mem[551] = 144'h04940454fb36fc6bf856fa88f611fcf0078d;
mem[552] = 144'hfb70f00f061bf4da0d14f08808d6fdf0f05e;
mem[553] = 144'h08c4008d033000c1f0fdf61f009404c7f755;
mem[554] = 144'hfad4087604a1f631f8e8fc72f0b0ff43f4c1;
mem[555] = 144'h0041f5d70b2ff06bf391f616f267082309c4;
mem[556] = 144'hf4e3fa060afc0259f08f06f1f99c0b8209f5;
mem[557] = 144'h0a5dfb1805af07cef164ff39ff75f3350e54;
mem[558] = 144'hfe50f3230b95fb01001cf5eb08bd08ed0783;
mem[559] = 144'hf335010f0ded08a4fb49f34c0080faaf0232;
mem[560] = 144'h0416f31709aa0d8dffcefd26082b0724f6c5;
mem[561] = 144'h0058062206fe0b0c05b808ff06f5f864f0f9;
mem[562] = 144'h07250337fa0ff2990f9403f5f7860357fa40;
mem[563] = 144'h0cd7f2ecf3bbfb74f562f88bf66401e4f861;
mem[564] = 144'h0cf5fcd7f356f880fbd3f31e0e9b0c2c073a;
mem[565] = 144'hf82b0a95f577f9e0f49bf9d0fa21ff5b0f35;
mem[566] = 144'hf7fffe62f293f9060f30fae2f698efd8ffd8;
mem[567] = 144'h0ff3f2b9f2f301a1f04df71005e003a6023a;
mem[568] = 144'hf5a1008d0e080b900f00f84a0b4503c20384;
mem[569] = 144'hf77708bdfb74001bf23dfe90f704f785f42e;
mem[570] = 144'hfb70f2f5fe77ffd5faff0d4ffb250037f0fd;
mem[571] = 144'hf606f960f8560d0df7770dd1f65af9f6f6be;
mem[572] = 144'h071dfa640c67f05ffa7d0a16ffdb01b5f7b7;
mem[573] = 144'h00f4f58bfdc1f3e9f07e07090c56094af079;
mem[574] = 144'hf284f011fe500b4cfd1708b8f9260cf6f5a3;
mem[575] = 144'h03f9f08f051bfe49054201fe00590685fcc7;
mem[576] = 144'hfc98f9f5f8a805040e490fc4f3b0fa61f584;
mem[577] = 144'h07f40337f2a9ff920b3bf1bc0079090af7b4;
mem[578] = 144'hf97c051c0f94059c0e3c0c5df93ef26b029d;
mem[579] = 144'hf7490aebfd64f6fcf706f9f0f741f24f02b6;
mem[580] = 144'hfc3604acfd4c00f201f9057f0991f9c8fccc;
mem[581] = 144'hf5a50834fab40f3cfc02f5f707a20a36fb06;
mem[582] = 144'hfe400f820cc2f4f50059fce4f50407bff40e;
mem[583] = 144'h04cb08950f9f0525fd5df2b2f883088e0620;
mem[584] = 144'hfbdafd540adafa64fdfbfebcfc1c087f07a3;
mem[585] = 144'h0d18f519f7ad0d6d0c08fedbf545f35bfa3c;
mem[586] = 144'h0b3c072c025ffc6d0d720559f5ff0d2df362;
mem[587] = 144'hfbc9f1a40444fcf4062df7470e08f6a00c53;
mem[588] = 144'hf32bf90c09c80db70ee007cb0179f869f5c0;
mem[589] = 144'h018103520cee089af09309da0009f37e0445;
mem[590] = 144'h056d09810b490abaf8abf8d7ef9402eb04a6;
mem[591] = 144'hf9fcfd92fa0c0ab1f13cf63204f0f6e20ec0;
mem[592] = 144'h03e5f84f0ae4f67a0bf8f6a8fb330e6df48d;
mem[593] = 144'h06bbf7e2ff9a01040b0806d6082ff543f3f3;
mem[594] = 144'hfb9ffbe9fa4beffff76b0f3df40bf0c5f59e;
mem[595] = 144'h0eeb057cf4ac0012fa7403930572f651f5e7;
mem[596] = 144'hf3d40147f7acf0d10aaefd21f50207420323;
mem[597] = 144'hf9fdf777fd8800a7f67bfbc90ceef15cf03c;
mem[598] = 144'hfb210314ff7c09b30c5c03890ce00c9df1da;
mem[599] = 144'hfc9cf5dbfe290454016907de04cf0cd30ad4;
mem[600] = 144'h03b8fe9b016ff6d10155fddaf0aaf8d704b1;
mem[601] = 144'h08b400e8fc47fe97001b079006a1f05c092a;
mem[602] = 144'hf42403bf0ed0f395f72bf6270998fd740c68;
mem[603] = 144'h0aa30f55f813f26cf5e000acffdbf711f3eb;
mem[604] = 144'h0c6c0166092cf661ff2af954fc790bdef48e;
mem[605] = 144'h0f170675ff65027b071308d9038ff68304eb;
mem[606] = 144'hf18df891f18ffad5037505c2f2b30377fa45;
mem[607] = 144'h06e8f98a097bf2860e650341fee4fccef488;
mem[608] = 144'hf8830d0cf24407c2f2d4fbd7fb8300450ec1;
mem[609] = 144'hf305ff34f682f7d70c1dfe5dfb4003f40783;
mem[610] = 144'h0d760b2cf757041b001b0176fab1fa2ff005;
mem[611] = 144'h0c42ffdb092807b7f10901410011f872fbe2;
mem[612] = 144'h099ff2e7ef7a0c110acdfc090dbbefeef1b4;
mem[613] = 144'hf762f72f04ff058f04aa0a97037bfbde0d49;
mem[614] = 144'h08c10a880c77f3ab06fef0480643016e0cc2;
mem[615] = 144'hf625f81cf0c90e54f0f8ff05ff28015afbb1;
mem[616] = 144'h0c09f978030ffa5901e203e4f42a0c9d0b96;
mem[617] = 144'hfe2104e7f5a6f038041f075d0059f81bf8fd;
mem[618] = 144'hf2780220066dfd4c0bd20ca60d48f2780353;
mem[619] = 144'hf141fffbf8d10d30f76cf2b7078300e80cac;
mem[620] = 144'hff9401a60d04f259f146eff2087ff3c0fdd2;
mem[621] = 144'h02baf85203080e540753ff5d07ad03b30086;
mem[622] = 144'hf6e4f7fe0d180a4702d9f0aefac8fad6039b;
mem[623] = 144'h0e1a095802b50947fe92f270f15c0462f89a;
mem[624] = 144'h04cf046701c006ef0e080151f36d01890bd7;
mem[625] = 144'h0d120bd4fbf604d80a3c09a7f26afa1afa99;
mem[626] = 144'hf699f533ffbdfcfe0a6a0353f552f8dbf711;
mem[627] = 144'hf745f42afcc90a03093f0f18045301a5f7f0;
mem[628] = 144'h037d0cbc0924f290fbd10f48f4170a6cf395;
mem[629] = 144'hf355f93502f3f641ff4a0b65f155fa740972;
mem[630] = 144'hf196f591fb6cf359f7b3fd03039e0f0ef299;
mem[631] = 144'h0d1a0abaf2d2ff0005710c380db70c170c75;
mem[632] = 144'h0a61fd4c0c4707900ed0fa9bf732f7e0fff9;
mem[633] = 144'h0bf3fad307e90b310598f37d01b002aa0264;
mem[634] = 144'h0caef623f9320bc6f6a9f3100fbff3110d7a;
mem[635] = 144'hfa200bacf4cff7130b1ef4a60320fa4afcdc;
mem[636] = 144'h04da03c7ff60f0ca0300faaf0bd8f3baff8d;
mem[637] = 144'h0d77f631035b016001c205b9fd42f2810131;
mem[638] = 144'hf52d09010c34f43a06900d91f910f3cc0b27;
mem[639] = 144'h0eb0044704e506320f5d02b304250430fabd;
mem[640] = 144'h0e56fc58fac7fc5c030bfbe8fa02067ff29d;
mem[641] = 144'hf21f016904df09fc023a0c360b73003200a7;
mem[642] = 144'hff35f81c015bfc66fc3004a7f5ddfba6fcf1;
mem[643] = 144'h07ed005805b40f120e640a82fd7bf885fc5f;
mem[644] = 144'hf422007a07f7fc8a08c6f79d0a54f274048a;
mem[645] = 144'hf1a2f3f4030dfde40e280473faea03b8f2a8;
mem[646] = 144'h0af3f5affc8b06c6f9d9fafd07abfbbdff8b;
mem[647] = 144'h0ac4f1830fcef76cf90af2fd059d076cf0e9;
mem[648] = 144'h00e00fd8f54e0dfe0e40f2d40ab20da9f02b;
mem[649] = 144'h05b4f9ab057af589f578f75defd207b5075f;
mem[650] = 144'h0f11fcbcf13cfef401dcfc77f945f1d30512;
mem[651] = 144'h0dca02e4ff5af6cb02760843f88ff583f7bc;
mem[652] = 144'hf550fce70793fd9c05010990f57a0e320bfe;
mem[653] = 144'hffd6f45cf6400999f9fffcbff2e6f5b0f766;
mem[654] = 144'h05ff02bef586055bf5abfb97fa13f2230a6e;
mem[655] = 144'h060f0fc9ff2bf6180655f340060df936fe38;
mem[656] = 144'h0baa0aabf1d503b70e01f2d9f7920253f596;
mem[657] = 144'hfadbf0d70eb20924ffb1023c0b220c2d0a97;
mem[658] = 144'hf7060cebfa1c08f1f62f06d7fe2c0299fa5e;
mem[659] = 144'h0ec003f50313efd4fa53f4dc085a09c9f32e;
mem[660] = 144'h065c029a0d6c0e7cf61f0b61ff900764fc22;
mem[661] = 144'hff680bbbf3370621011c08b2f4def377f220;
mem[662] = 144'h06b2043e02d2013d079e0dc3f5d10dfdfa5c;
mem[663] = 144'h0510f5a506a707bb07d80329f97f0be203e5;
mem[664] = 144'hf87c0a94024e0238f7a00d8cf1bf0782043d;
mem[665] = 144'hffdf0e11f33104d30da802dbff58f050fad7;
mem[666] = 144'hf2800d3f04d00ecaf87d0bba0277ff53f58f;
mem[667] = 144'h05570eb60a92fafafbe90da604e2ffe0fa51;
mem[668] = 144'h07b509a00dce042301790e0df00e069d02c9;
mem[669] = 144'h05610eb90fb0f995fdcdfc4cf54c04cdffc1;
mem[670] = 144'h0808f3d50d05fd910ea0f4160e22f2d3f1ff;
mem[671] = 144'hfc330175ffdaf9c0048dfd97f22afb850a86;
mem[672] = 144'h05a3ffa0f906f17a06d1fcc6029304f9f9bf;
mem[673] = 144'hf2a709e5ffef018dfb720d0c0f790d820c04;
mem[674] = 144'hf345f60201af0f61fe99f01c0c54001c005f;
mem[675] = 144'hf80ef17ef0dbefe5f3f2ff05f2f70d42029a;
mem[676] = 144'h09df0e100bec0b17f5b00a7d03a6fe06fb7a;
mem[677] = 144'hf1250d9cf904062b02f2fd74fe150088fc0b;
mem[678] = 144'h0924f76e010b0d460c5c0a9c07a105a30a04;
mem[679] = 144'h0caffff50475fa4bf53c05e90496f9110c85;
mem[680] = 144'h0088ff70f7f1f1ad0acdf3fc0cd6f57b0f29;
mem[681] = 144'hf4f204bbf8d80eb10fd7fe57fe4ef203f446;
mem[682] = 144'h0143f80ef30803edf2e1f01001e102310c3d;
mem[683] = 144'h02bc0a2600b80e39048c0ac6f3a6f878037a;
mem[684] = 144'h04c2effc05fff7fd0068fd23f53eef5d059b;
mem[685] = 144'hf426fa20fd25082a0bd6f89d02f1fbf1f8c3;
mem[686] = 144'hfeb40c7cf1c2f2f000bbf693ff57fa5203bd;
mem[687] = 144'h04f10b450192f17c02dc0f1e0d59f321fea4;
mem[688] = 144'h0a070ab9031bf8770c0204d60e3e0c84052d;
mem[689] = 144'hfa83f94df7f90848f96bf0b1f04603a90032;
mem[690] = 144'hf900fe1101c206aa0e090dbc0dd50132f86a;
mem[691] = 144'h08010a0ff289ff9f05b7f621f24ff5a10fba;
mem[692] = 144'h0877f2b5fe7e078e0d86fee9f82701ddf168;
mem[693] = 144'h03c7f1a6066ef9430f430fa60b2df5e8fe16;
mem[694] = 144'h0923f14806e10e1dfa950285fbb20636f703;
mem[695] = 144'hf3c706cb0ccd061cff350aa5f718f97a02f0;
mem[696] = 144'h09cafaf1f4bef584fd97f9d5fde9fd85041f;
mem[697] = 144'h0532f4b7f58308edf097f2530398fc10f0e4;
mem[698] = 144'hf38108380908f847fc60f0faf28ff3e3f0ec;
mem[699] = 144'h0d96f42bf5a7fa150c9dfd4201c80722ffd5;
mem[700] = 144'hf28903050fd7fce7fa76fa78f997fa91f7ad;
mem[701] = 144'h06430f3d0915f20afdd60e13f4f7fba3fd3e;
mem[702] = 144'h0b1ffbb10315f013f4d30ef10524f83cf630;
mem[703] = 144'h06780355ff6ef93f0002fb5b0d8af1f4f48f;
mem[704] = 144'h0383f38d0445f39605fd02dd01ab01b907ef;
mem[705] = 144'h0fde05ecf5f7f3890553f993fa5bfd0705e7;
mem[706] = 144'h072e07eb02fa04bb08ef0f20f3c3f1760488;
mem[707] = 144'h01fb09ddf0220822fd6ffea3f5f40a39f4d3;
mem[708] = 144'hf11d069cf864f37bfdf4f7cd08710a10f41e;
mem[709] = 144'h07d6f3810e5806b100830afa007702a7f6bb;
mem[710] = 144'hff30f0740f09fb0302d2f8edfea60d900470;
mem[711] = 144'h0188f04104a1f839f157f64cfa6d09800ab2;
mem[712] = 144'h004cfaaf00f3f19e0c99f2a60910040efa65;
mem[713] = 144'h009ef1330e28f9faf400f59ff2bdf0cb02b3;
mem[714] = 144'hfd470bda0057048ff296051bfea0f7d107ac;
mem[715] = 144'hf5a4f6de0c45fbeff2f4f8080eb4f245fc84;
mem[716] = 144'h02fe0839054afcb1f42500160bf9f4860cee;
mem[717] = 144'hf9fcf6b5f27af1320a28f1c1faef0199f69f;
mem[718] = 144'hf0020235f6540d82f3b0fdc8fc96f27dfbc7;
mem[719] = 144'h03c500320f6804fa0896f5c10ff202f00f48;
mem[720] = 144'hf87c055b0f0f0f7bf293f276fc78f80ff36a;
mem[721] = 144'hf60e0654f41dfc3d0cd1f7f80b57ff050e60;
mem[722] = 144'h0884f9ae04b6fae0fba40eb4f1a40eda00cd;
mem[723] = 144'h0fadfa290196fb13f2e0f78607a1f739f725;
mem[724] = 144'h0d450048f46008f203f0fd0c05fff4d70157;
mem[725] = 144'hfd14f6730c74fe9af05ffbab0b5df0030811;
mem[726] = 144'hfd86f72bf38ff9190d02fd87f6edf4a4f623;
mem[727] = 144'hf9f8f67405c8f2cc029cf9fefc9404260b1e;
mem[728] = 144'h09fe0ef50f6404d1f053f716fdcc03f40bed;
mem[729] = 144'hf2a80af2f6fe0675ff4d034cfc8ffc85f292;
mem[730] = 144'h09ad0b35f1e607d1f52c08deff320b500c25;
mem[731] = 144'h0f700aab0c5ff6210267023905d8f634fbf6;
mem[732] = 144'hf9b70803f79c05b7016e0526f43e028cf0f0;
mem[733] = 144'h0478f17cf7780eb7fab0f424fde80b24fe2e;
mem[734] = 144'hf7b80539fb3004adf054fc81f2b505ea010b;
mem[735] = 144'hf74bf8ecf762fdfbf525fc97029a0294f85e;
mem[736] = 144'h05ae03390333fa6bfebff0670d450515f1ba;
mem[737] = 144'h05eaf71f09cf026e07f9f8aafd8afe6e0cf2;
mem[738] = 144'hf56702c6fd9a0d5cfb34fcba010d0df70096;
mem[739] = 144'hfb7ceff4fffd0b91097f04810e88f5630722;
mem[740] = 144'hfaed0431031d05720d6907f9efc707160acf;
mem[741] = 144'hf2f5009afbaf0249f88e086b0d5f0f25f598;
mem[742] = 144'h0dd4fabff69b0ee1f1d1fb8508a1f0a907ce;
mem[743] = 144'hf33801aefc73f9f0097f0bc1059ef5e8feea;
mem[744] = 144'hfc760d3b05fb0ed706260c940f58046504b0;
mem[745] = 144'h027a0e42f9b2ff7600580aa7f31afa630d21;
mem[746] = 144'hf3380dd2f4c80e05f6b8fdfb0875f26104b3;
mem[747] = 144'hf231feb609620339f12807ff0718021e04ff;
mem[748] = 144'h0b5c04a30845f199feb500e2f7e50692f52e;
mem[749] = 144'hf17f037d006d0b6efaf8072ffa66fcfef314;
mem[750] = 144'hffed0724070200fd08b3043efef600320c56;
mem[751] = 144'h0e06f90d0e190819f102f9e6067bf535f648;
mem[752] = 144'h0e9f08aaf9bf06ed0e98074afc08f5a8efda;
mem[753] = 144'hf63efba8fa97f0900ba70127ff3105b1fb00;
mem[754] = 144'h013202750aa40105f11807540bcff1a4fc8a;
mem[755] = 144'hf8a60331093f08c504aa0a160032070c03a0;
mem[756] = 144'h0bfd0ea008f8f828f985f1690b7bf5270b65;
mem[757] = 144'hf5c505ca022df82effa001d7f2d6ff4bf76a;
mem[758] = 144'h04b6046f00bb0d2002b307020e3e0e78f631;
mem[759] = 144'hf23900a60982fe7af076f717fdaaf653f1d3;
mem[760] = 144'h0a7ef315f4f6f18bf6a90be6ff4cf7520a22;
mem[761] = 144'h08530186f15ef296ffa90cc9051afe8af409;
mem[762] = 144'hf16bf7b00cd30f860e5ff2990e2503e3fc18;
mem[763] = 144'h0ce50ec207140cee0c8a06b70d16fe6af5fb;
mem[764] = 144'h0facf8d8f9620c2df6f504a60188f127037a;
mem[765] = 144'hfbbe0b3900090dcaf8340b740c8ff548f21c;
mem[766] = 144'h0236f8920702faff04950b080cd7f8fbf76b;
mem[767] = 144'h0826f4c10ca8ff32faf3fa4cf8c204460e18;
mem[768] = 144'hf738fa27f59ef83c0ee80871f1f9fcd3020d;
mem[769] = 144'hfd70f18a0e170632f5d4f3010e7606b20bf0;
mem[770] = 144'h0f23fdb20c71043f06f6070a0210fd110f24;
mem[771] = 144'hfad207100eca0b4cf7f2f853f1010445fb3d;
mem[772] = 144'hfc9e0d47f28cfec501d0fbc303400ecdf059;
mem[773] = 144'hf29f035e08ecf84afb7500c80fb6f59f02ab;
mem[774] = 144'hf822fb1df989063ff06b0acdf6ec0c8ffd55;
mem[775] = 144'h06bcf15cfd320ddcf20d0a56f2e707e804c8;
mem[776] = 144'h0508f70fffba057ef97a0f91fbf70d1eee76;
mem[777] = 144'hf654ff28f759fc58fc870428f1e800c90e93;
mem[778] = 144'hf4b3f35e0562f4530a010bb806b4099701b9;
mem[779] = 144'h0909f7b60cebfa560a1af59600de01b20187;
mem[780] = 144'h031afec8fd4df676f68e08b7effff51cef20;
mem[781] = 144'h02be0a2a04a9073bf070fb4a06b3055bf23f;
mem[782] = 144'h00bef06cef4406130b75fe5ffbb1f3df02fb;
mem[783] = 144'h0e9cf061fab508a80a7b00630f49f90d09bd;
mem[784] = 144'hfed70a11fbb9f752f970f9710401faf40b12;
mem[785] = 144'hfa9206b1f4090b4b05ee0380fd4003e0f300;
mem[786] = 144'hf0580e14f37ff262014af37e02810684f166;
mem[787] = 144'h0038fcf70d40f1adf1e600f7fa7105250ff2;
mem[788] = 144'h053cf4f4f9ebf6b40d15015ff286f506f41c;
mem[789] = 144'h02e2f018fe6807c5013f0c110551f83803ae;
mem[790] = 144'h0d49f039042b0233f01af0dcfdb3f7bdf12e;
mem[791] = 144'h0ecb0912fc8df4b5fef1fab601380dba0319;
mem[792] = 144'hf390013af24ff09bfeb906640bfdf693f688;
mem[793] = 144'h0220083e0cf1f2b8f2cdf94cf80b0654f039;
mem[794] = 144'h033f00540b56fa21fddb0e8afb320a7df294;
mem[795] = 144'hf9fc0d2df6a704fe07b5f9fefb77f855fa38;
mem[796] = 144'h0b670c9bf1a3fce9f06c0528f2c507d008db;
mem[797] = 144'h07e4fec1fff4f25a0f2d0f750c6405c0fbd9;
mem[798] = 144'h025100bef2ae014f0e3cf7e0f6d207ed0688;
mem[799] = 144'hfed70970fda50c12fc8bfeaff1d80ae30664;
mem[800] = 144'hffef09970513f41cf2fff019f46e07f5f1b9;
mem[801] = 144'h08e2f59502e9f30303c605140033f016fc46;
mem[802] = 144'h0f010854f9c8fcb0f652f6290a8009c2f204;
mem[803] = 144'h0be5fb3006460e7c0730fb5c005b06cdfff8;
mem[804] = 144'hfd9a0b4a013ffb7c0d10055bfd47f525f83a;
mem[805] = 144'h094207b1fcf7f43dff840aabfa31efe00846;
mem[806] = 144'hf3abf63a086807effeaf040402de049706f6;
mem[807] = 144'h073906ab0e7b0a0df6b2fcd8fc7af0420667;
mem[808] = 144'hf5310e39fa720e6bf71df385fb3cf8fb0a61;
mem[809] = 144'h098ff337f728f1be0eeff774f15df5d00a3e;
mem[810] = 144'h087df918f9a3f86609670eb1f4760c2ff215;
mem[811] = 144'hf45200b0f93907440f8ff2c3010cfeecfe0e;
mem[812] = 144'h00b7fea4fd5ff99ef5f40c99fe020461fb77;
mem[813] = 144'hf956059509a70e94fcc90c9501c1042bf785;
mem[814] = 144'hfa35f70bf87b0708041f066af4a408450c74;
mem[815] = 144'h0fa0ff8c0735f1a5f5600692fbaaf5cbf626;
mem[816] = 144'h0d1a0b65fdae018e0c81049e0a20f65cf948;
mem[817] = 144'h0e4e05b40eaf014a0636fd370e25f725ff4d;
mem[818] = 144'h081001ee0f0f0a090390fb6afd00f993f98f;
mem[819] = 144'hf0e40a81f566f13f07ebfea2f96ff27205a0;
mem[820] = 144'hfcfffd2bff4bf0b4fbcbffc00d8df27d085e;
mem[821] = 144'h044801e5f449f323f950087ffa45f56d0e50;
mem[822] = 144'hf60b0f10fbd3f67200cd0983f12e026ff296;
mem[823] = 144'hfbc80611fde10a1cf1db08a4025ff7b5016d;
mem[824] = 144'h084a0aa705b9065007b2f9110844fc230b9f;
mem[825] = 144'h0e2ef8a9f7ab0a440d3907c90b7b0c0c0855;
mem[826] = 144'hf315f04af252fedcffc4f7a8fc4908dd0265;
mem[827] = 144'hf4570c6efc390d0af55f05fe080cf1c8f16f;
mem[828] = 144'hf8afffec0c39fa10fbf303c7f7aef087f1cd;
mem[829] = 144'hef54f5c7095c02630774046c06f5f55d0036;
mem[830] = 144'hf1c6f515f286f5ecf8a5f3a409770c1cfe81;
mem[831] = 144'hf0cc091ffedbfad8f026feceff2f0c0e048b;
mem[832] = 144'hf153f81b036c02960199015907e600f20d92;
mem[833] = 144'h04e6fb5efc1bfc99fd65f3b00f0f019304c1;
mem[834] = 144'hf78af145061d06d6f0a2fec6f511f59601eb;
mem[835] = 144'hf3730f2e06460575f274093dfe3affeff4de;
mem[836] = 144'hf751f038fd3905ef0d71f8f1ffc30ed5f2e3;
mem[837] = 144'hfc49f321096807560c850d8b09b1f0b9fbdc;
mem[838] = 144'h0a30f248fb530884f0fe02d809120c240e3e;
mem[839] = 144'h078ff0d90dba0d9ff0c2f4000f1af0d4f161;
mem[840] = 144'hf6b8f36a05df046d05e9f4f8f50efd0409e5;
mem[841] = 144'hfe990bcef936f4f305bc0075fd71fe9f0bb8;
mem[842] = 144'h08e70a8afac2f0aefa07fc35f2d9f72204b5;
mem[843] = 144'hfd05f6e70474f0f9f9cff85705e60cad0e1e;
mem[844] = 144'h0824072102db0496ef6801b1fc3d04f1fe48;
mem[845] = 144'h0f00f313f8480281efcff52601da0f40f700;
mem[846] = 144'hfc8bf299f5fbfca7f145f20df52a045e0835;
mem[847] = 144'hf0d60554f8b6f5acfb3c0d440465fbd4f0e6;
mem[848] = 144'h008df04b08daf402f2f2f92df0430ddff910;
mem[849] = 144'hfddb07e7f5caf1ecf2680edd0aa0f104efb9;
mem[850] = 144'h00710a19094907d7faf10b6bfc55fd4cf79c;
mem[851] = 144'hf1800ca6f2b404da046e00a8f43a0d56090a;
mem[852] = 144'hf1b4076b070ef2ce0271fdfff7a90ef60023;
mem[853] = 144'hf07cf2c1fffa0b6a06cd0db90b89f0f80f7c;
mem[854] = 144'h0c3ff1b6ff8b023a021def4304f50e79fc9c;
mem[855] = 144'h0dfefdfa00d9f45d0386f896059c052ff380;
mem[856] = 144'hf4670a140b8900380a2df15d084108470025;
mem[857] = 144'h0da7003dfd470889fb770c820cbc0cabf6fa;
mem[858] = 144'h0722f859f50100c40ae808130791030ffd46;
mem[859] = 144'hfaa9f58ef7d0f23cfc9b07ff030a0d6ff559;
mem[860] = 144'hf0d2fab00b1ff7d8f01ffaa4fecbfed00af2;
mem[861] = 144'hf54901cb00ea0645f933f0ba0d70f17f08fc;
mem[862] = 144'hf168f2150590f43b0cb60ca7fe01f33ef562;
mem[863] = 144'hfad3fdd1f3b1f96dffabfb01f71b0196f860;
mem[864] = 144'h068b0a2cf836eed50350034e0c0cf7e0fc44;
mem[865] = 144'hffb9f8ec096ff1c70b0b03b3ffe90ef9f5a3;
mem[866] = 144'h05e50295f1a7f923f1a2f1a5fe66f159f8e7;
mem[867] = 144'h01b406d3010b0359f2ad08d305afff0e0bc2;
mem[868] = 144'hf740ffc7085c0ba308f50dea0fa20d85f4f2;
mem[869] = 144'hf79f09b8fd66fc51f1110ce4f864f2170564;
mem[870] = 144'h0967f28001abfb42f4910034f0ef0c16015b;
mem[871] = 144'hfa4904d5063e069b0502f1fdf95302910e09;
mem[872] = 144'hf6f303700f51f1f5fd4df556f21ff60df7ea;
mem[873] = 144'hf980f500f66b0571f0c9faf40246fca80b9f;
mem[874] = 144'h0f4106a907c9f18a0296f40bfe9bf135f193;
mem[875] = 144'hfcd2fe39f20c0ab603c702b70ba4f47c041f;
mem[876] = 144'hf6960bcb0b490e820aba0526fe990a1fef45;
mem[877] = 144'hfa06f182f55dfe4209700c63f5ae05760079;
mem[878] = 144'h0d2bf274f774feed0890f02af197f5a10f51;
mem[879] = 144'hf7960caaf13bfaa3fe080730fdb7fe19f910;
mem[880] = 144'hf20affcaf83d066af321f36cf8fceef4f51c;
mem[881] = 144'hf5f807d60887f746f41d000402d8018dfdda;
mem[882] = 144'h0630f2290751f4b405080f0a0e0ef4fb0a9c;
mem[883] = 144'hff4a02e40ee3025a06c605f20985f678f4ff;
mem[884] = 144'h0f1dfd430aba0a5af774fcf0f32601cbf553;
mem[885] = 144'hfc6509bef578fd27055ff7da0b050501f3f2;
mem[886] = 144'hfb04069d01e10484f322f5ec01b105f7fbc2;
mem[887] = 144'h0289034ef285f4c1f432f9380382f6d5f0c0;
mem[888] = 144'h0e000e1e0902ff2d02b306a5f52006720ac2;
mem[889] = 144'h0bfbf5e7f260f47503f7ff37f2410fb60df6;
mem[890] = 144'h03bff31f09d2f047f54702cff4c6045ff15d;
mem[891] = 144'hf40002e204c90caa0895011909d00076fb9c;
mem[892] = 144'h0aa4f6670d2cfff6f258fab7f5180cd2015f;
mem[893] = 144'hf715fd3107c1faeff07bf22d0b4af1c9067a;
mem[894] = 144'h02b8f7f2fae903c3f78bf8390c26f3ccf6d0;
mem[895] = 144'h021505cdf4a0f8b7057a06e2f208f11500e7;
mem[896] = 144'h090a006efb3ffe6ef141092e01eaffc1fafc;
mem[897] = 144'h029b08ac061bfec0f307058c06d00c4d014a;
mem[898] = 144'hf87cfd6ff49ff3abfd7cf8310c7cf763fb8c;
mem[899] = 144'hf474efe0070bf8e808db0b340dfdf2aaf3dc;
mem[900] = 144'h0724f7a90bec0c070304035bf995fe14f0d8;
mem[901] = 144'h0d56f14bf7f705bdf9e6f5d60c76067afec9;
mem[902] = 144'hf173f39709b40a89fcae0b40fbeff5fc0f4d;
mem[903] = 144'h0e1800e1f987fa42040c09abfd61f7fd0a73;
mem[904] = 144'hf7a7f43c04f10d53f03aff4e07b7fca6ff38;
mem[905] = 144'h0270fc5e0f44f4f503910b520967fe68f161;
mem[906] = 144'hfa7e074808c103b0f8990d32f0bcfdc30ce5;
mem[907] = 144'h0052012e08c70c71057201b20359072d0ff1;
mem[908] = 144'h05f10aed0553f8fcfafe095d0c7f025af812;
mem[909] = 144'h06160f470c7ff599fc87029ff912fe6cfa76;
mem[910] = 144'hf48007eff445fcb20093f526f8abfad7f286;
mem[911] = 144'h0e7ff670f06a030a0850009df554030102b0;
mem[912] = 144'hf61eff750b41fc92fedd052b048005220c6a;
mem[913] = 144'hf2ad083c0be60ba30b5300760d3d0ea5ff58;
mem[914] = 144'h07d5025ff1570379f253f399027cf1ec06f4;
mem[915] = 144'h0248f847ff3a0f270e17f15f07000d4cf45e;
mem[916] = 144'h08060bf20d4a0bd90538f656f4dbfffbfe54;
mem[917] = 144'h0cd9f1f4083bf2ab074b0949f5a2030cf298;
mem[918] = 144'hfa0ff7d5026e02490e7f0981fc67f36ff4b9;
mem[919] = 144'hf19bf2180cb00b58f698061301c5f353000d;
mem[920] = 144'hfa6d00220455f41808060daa055afdcffc0a;
mem[921] = 144'h01f5f419f11efbe4fb2603370ba3f4ebfd64;
mem[922] = 144'h0bec0445fe4c0789f72b056cfd22fe3df675;
mem[923] = 144'h0edeff5a016a0a06f8520889012af47c03d4;
mem[924] = 144'hfaec07f50b6cf65b00ff0352fcfd0b83fa2c;
mem[925] = 144'hf98cfdc60c3efa400eedf57c02e104410978;
mem[926] = 144'h06c8f955f485027bf234023c0c31fa16fa70;
mem[927] = 144'h0a17f7fff58ef60e068bf3bb00d8f9e709ff;
mem[928] = 144'heffef9e2fff4011d043bf6ea00fef61c0d37;
mem[929] = 144'h082ffbc0ffbbffce0bbc05210f7ef70af4ff;
mem[930] = 144'h022ff93dff5cfb38f8530fc1f4b40d83ef97;
mem[931] = 144'hf81afae70084f3cdf92df9d6fc08ef3504f5;
mem[932] = 144'hf417f69908ea00ef04bbf1d50c06046c0949;
mem[933] = 144'h0d49fce2fbba00da0c6906e3f470011df31a;
mem[934] = 144'hfab0fdf6f861fc78fb09ef5f0b1b06320c08;
mem[935] = 144'hf763088c0bb608d0f5f8ef06f02001cfff73;
mem[936] = 144'h02a90bc908ecf12806ab03b40717099c092d;
mem[937] = 144'hfa420c6f0e7bfa67fed7f970ff24f6e8f62b;
mem[938] = 144'hf3350db0022bf4edfef10a760b0c00b3f0f8;
mem[939] = 144'h0f5bfa4cf36a034302290aa80821f98cfd5f;
mem[940] = 144'h07ccf094f5d3f73b0aaa0204fc57f36ff56a;
mem[941] = 144'hf33e05dffaa8f051fbde0c210c0cf1d6fef2;
mem[942] = 144'h0a8d09ee02f7f7490c3cf81bfa13f9c8fd5d;
mem[943] = 144'hfca6f676037ef414fdc1fddef11afaf20b8e;
mem[944] = 144'hf7400010003f06db06d1f1f2093af4b5f5ad;
mem[945] = 144'h0f430d0cf3fd06d9ffa0075b09130535ff16;
mem[946] = 144'hfa8908a0fb4e0e11f89cf636f96306c3fb35;
mem[947] = 144'h0f04f62cf47b0c07f9320656027eff77f808;
mem[948] = 144'h0e1ef9f001410dce03d0f41f0622f36f057f;
mem[949] = 144'h01d4fa090969f97dfd2e0c8ef659f1faf469;
mem[950] = 144'hf81d04f00d2909fb002cfa16078e0177f414;
mem[951] = 144'h0ec404b8f5730fa0f6090715fdacf3fff276;
mem[952] = 144'h01030d9efec4f46806cefa200b6e0134020a;
mem[953] = 144'h0eb50e320ab8ef5701caf089f2cef28301f2;
mem[954] = 144'hfab00ad80705f30c0b95f14002e3f99501db;
mem[955] = 144'hf05e0ea1f8c00f8afe400ee50389fc6d0257;
mem[956] = 144'h094601da0beb0179f620fe060d9c031a066e;
mem[957] = 144'h0b6800fe0bbb05300e33f22ef441f3980133;
mem[958] = 144'h08a7fc720df00ba3f57d0cb4f15cfc0af603;
mem[959] = 144'h0859f6620dbe05dbfa2e0c76ffa2fa5701b7;
mem[960] = 144'h0180ff7b0ef2016bf31d08c50da4020a0b4b;
mem[961] = 144'h01c00e3d01db0512f4d7f1c4f40606bcfa8c;
mem[962] = 144'hfaea0dc3fd2d01e7f0f3f9ff042df755fa54;
mem[963] = 144'hf0d9f7d801adf13303c90ed607ad08ad01aa;
mem[964] = 144'h0c47fbe2f00008160348f08cfef5f5da0d1f;
mem[965] = 144'h08ac0345fbee04c6fa2dfc52f5ddf5510501;
mem[966] = 144'h0f2bf87d06e10a2ef4cf07dbfa9c0419f17a;
mem[967] = 144'hf76df21af74f0d940556059d0743fb6503f2;
mem[968] = 144'hfca4077c0eddf292f90bfaef030b0333f8b7;
mem[969] = 144'h0c28f787f92ffb01049ef604f288f72bf062;
mem[970] = 144'h04affd48fa0df6c903bf0dfbf550062dfef7;
mem[971] = 144'hff1ff9a908990bac02ce04ff089ffaff0b73;
mem[972] = 144'hfc820894fa370698efe2fe71f3b3f164f3ea;
mem[973] = 144'hf538f42104a8efff0a0f0e77018cfc9af799;
mem[974] = 144'h08dafc3efd74fe83fa95f01af47c02130655;
mem[975] = 144'hf993030307e7080a05de06e90d91fb1901a9;
mem[976] = 144'h0f89f57b0514f827072a024e064afd1bf771;
mem[977] = 144'hf4bff334ff6af699f543f3cf0d1bfa32f886;
mem[978] = 144'hf93d09f80e230b17fdf309860d11027af8f4;
mem[979] = 144'h018f0786ffcafce20bf40e090530064df3cc;
mem[980] = 144'h0d50fbf90f5106c6f281f9c1f4e1036f0c33;
mem[981] = 144'h093ef7ef0858f0c7f887fc14075ef737fe50;
mem[982] = 144'hfd68f606f4ecfad3f98f02610807f826fcfc;
mem[983] = 144'hf9a6093dfe95053f08ad0be5fcef03bbf208;
mem[984] = 144'h0f87fcb9f9b3f8ae05170511040ef92a0230;
mem[985] = 144'hf91ff9d303dbf8c8095af80009baf7b6031c;
mem[986] = 144'h08cefef308e7f3210755f53007660ad5f82c;
mem[987] = 144'h0dd8f105016800dff18cf38bfffefd86f3d9;
mem[988] = 144'hfd68ffdf0b6e0f61f62b01f8f4fc0c6c0c26;
mem[989] = 144'hf66ffb02f434fcb0f3d9fe2f0cbeff52097a;
mem[990] = 144'h0365f9f405d2f59eff13f79505bef904f2a1;
mem[991] = 144'hf0db08c40f510fe20367fe15fa32f4f3fe0c;
mem[992] = 144'hf11a019bf4320c62ff5afa8609cbf98f0074;
mem[993] = 144'hf1cb073e0f480f2f034a0cc2f15df983fdff;
mem[994] = 144'h0585017b0ba4f79ff438fac405daf4c80d60;
mem[995] = 144'hf5c2f8f0f8a60a210c120530fb98fae70d20;
mem[996] = 144'hf093feef0cb9f5d1ffc7f36efb4f0a1e0121;
mem[997] = 144'hf57ffe8d0376f9c2fb94f903f274f42cff63;
mem[998] = 144'h060f0a7503f1f2c60c11f34f04ec0bb2f3d0;
mem[999] = 144'h0851fda302d1febb0a12f1370edefac80bcd;
mem[1000] = 144'h00a6f2bafbb7fa53f4ddf2d3f0c1fee10c41;
mem[1001] = 144'h0dd20f28f376f885fd7efe600050f0210b14;
mem[1002] = 144'hf69bfa24fa05fb9c0a77f32df94e0de5f3ce;
mem[1003] = 144'hf00e0862fa5eefec0188f41d062ff71d06a2;
mem[1004] = 144'h004c0ec309d1042f0ad4018bfa9209240b08;
mem[1005] = 144'hfb8cf0060dc3f05a0bc10e26015df5150941;
mem[1006] = 144'hf23e09ad03c4fb58f708f1e3057300a105cb;
mem[1007] = 144'h054801dbfdb4ffbf087a0956fbb7fa2b05b6;
mem[1008] = 144'h01b5f6ebf90afdc30bba0271f97f0a99f349;
mem[1009] = 144'hfcc90f44037c0c950d3d002406e0fb8df4fd;
mem[1010] = 144'hf0b6048cfa8309d50da80128f6e2f0cff95f;
mem[1011] = 144'h0a600a1bf6f4046ffd08efd6f121f5e10712;
mem[1012] = 144'hfdbc029af9e60629f735051907eafccbfcb7;
mem[1013] = 144'hfac1fc2cfef3f41f0f1dfbc70c5cf4360f06;
mem[1014] = 144'h0edbffe8f4e1f5fa06ff06660648f3d1f29f;
mem[1015] = 144'hf919f44dffb10051ef8ef40607aa03e2fd82;
mem[1016] = 144'h037703c5f5f90007018d0971fe94040f02cf;
mem[1017] = 144'h0d2df7ca03f5f5110189fbcafe4808810283;
mem[1018] = 144'h0d6c0923f7ce0d06f0090e910800f771fd43;
mem[1019] = 144'h086efecb00830e92fed904bf092f02de0045;
mem[1020] = 144'hf4c9faeefce80d510e10fa80f4e9f257eff1;
mem[1021] = 144'hf1de0edaf35706e206280b97f165fa5bf66e;
mem[1022] = 144'h041a0630faf2f9970bec00a106580443f88d;
mem[1023] = 144'hfc710825feb00afdfffff95003dffaa1fa61;
mem[1024] = 144'h0cb7089203e50cb1031cfe1efb02f4810689;
mem[1025] = 144'h0cb1f9d00d69fe82ff55f25c0f9300fe01b0;
mem[1026] = 144'hfd0af36b02d5f883f4ff0095f6e70643ffe9;
mem[1027] = 144'hf895f44400cbfc39f05af27efb6c03f3050a;
mem[1028] = 144'hf08103ba0182075cf076f26ff6ee03aff385;
mem[1029] = 144'hfc0401a3fd5ff844fe69f7a0f3f90d73050f;
mem[1030] = 144'hf36f010ef761ff8202390cba0e650ca3f568;
mem[1031] = 144'hf85402f60ccd004c006a0b7501cef147f24c;
mem[1032] = 144'hf33f032af3f8f2b6f6c9fe37fa3df80d05e5;
mem[1033] = 144'h0d670aae0a74f8e9f178fd740b00fefaf753;
mem[1034] = 144'h080d036ff8980013f253fa9fface022ef825;
mem[1035] = 144'h05800d2ff80a0ea10c6d01ed01ca090b0b0f;
mem[1036] = 144'h06080bc20adbfddc0989fc42fe04f3d903dc;
mem[1037] = 144'h0949f01101fff94bf7780e010d050ce5ff13;
mem[1038] = 144'h029d0219f4e704d006530d6f0dfc03eff5df;
mem[1039] = 144'h0cd904650f08028a0670f2dcf7580c320c71;
mem[1040] = 144'hfed701f7f7eb0a8ff2ccfafc0afe0d0607a1;
mem[1041] = 144'hf8620c4f01390c9c00eb04af042809620a52;
mem[1042] = 144'hf0110f970501090903b30bbe0336f87cffc7;
mem[1043] = 144'h0ef3ff970128f420fc30019103bafd02f56b;
mem[1044] = 144'h0dba01e6ef7bfc870d8eff04fe45fdb102c4;
mem[1045] = 144'hf5bf0223f9d8fb1a0a69fdb1f391fc10009f;
mem[1046] = 144'h021bf90305b805e808cb044b0bcef04c025c;
mem[1047] = 144'hfcaafa9806900c6ff0be08650066fef2f700;
mem[1048] = 144'hf0f9075705e1fde7f25dfbb5f3af048d0cb5;
mem[1049] = 144'hf61304d00b86fb15efe4f9a0067c09360c65;
mem[1050] = 144'hf89e04d0f89bef77f4160eec0b7af64d0740;
mem[1051] = 144'hfa580544004508b6062a025a00d0f7bbfb22;
mem[1052] = 144'h092903820a110a96f9fb065cfac40bb60197;
mem[1053] = 144'h0388f85600460865f9a30af4f83a0078ff78;
mem[1054] = 144'h07dcfd35fe36fe3ef943f7d1f3ca087a06df;
mem[1055] = 144'h0fdd02ea02350af9f3baf980020603a30e5b;
mem[1056] = 144'h04db0aecf76afaee040c0c800522f58f02c2;
mem[1057] = 144'h08d30f54f7f7feba00c2f55cf398066e0aa9;
mem[1058] = 144'h0be0fa7c01f9f8d405affc3909b4f7100d3d;
mem[1059] = 144'h0cb00f62f3d0fe7bf6ee00a5f57f017202df;
mem[1060] = 144'hf5640d8ffa84fc87f38100d30900070b0f5f;
mem[1061] = 144'hf0ad05aaf0dafc4f0d63f9e0f5d70e370c17;
mem[1062] = 144'hfbfefd6d0f3a05010f6d05c2f696f51f00ad;
mem[1063] = 144'hf8700f5908e3074a0fd508dff380004cf049;
mem[1064] = 144'hf3650137f0590c3c016e06a2f741fce90be1;
mem[1065] = 144'h0b57f069fd380e4df4160894f65608c6ffbe;
mem[1066] = 144'hf93b0a7ffd3bf6db0453f099fec0019d0cef;
mem[1067] = 144'hf98e0f38f32105acf9a60588f9830538fde8;
mem[1068] = 144'hf4c70c33f27d0a6107adef9bfba300cb0ac9;
mem[1069] = 144'hefbb07ea0194ff5bfb030b0af0e5f1a20cec;
mem[1070] = 144'hff11f056f462fec0044807a503b003580919;
mem[1071] = 144'hfcf90a42f44afba4f96109f80533f32bfdc3;
mem[1072] = 144'h0879f35bffdb0bd2fae2fb230c3d0b82f7f4;
mem[1073] = 144'h08260faff3a802cff1d40cc309ea0a69f299;
mem[1074] = 144'hf76809e90533f5c4fc29f6a3f45af34ef729;
mem[1075] = 144'hf6f9f5affc070ec304250db8faa20ae7094b;
mem[1076] = 144'h0138013df8e806f7055af3f0f9fd081dfb37;
mem[1077] = 144'h0c52f1e2fc74f4b4059208400b4afd65f7ac;
mem[1078] = 144'h0e0cfa8f005cff81f01c0498fc7006a2003a;
mem[1079] = 144'hfd6ff5af05ef01be0803029d0b530a60f936;
mem[1080] = 144'hf057096b00c0f54e065ef91a0adffbea0881;
mem[1081] = 144'h031af541f8250ebf0fb2fdeefb7efb620c66;
mem[1082] = 144'hff6ff446fd47f82ff9edfe0004e304050c99;
mem[1083] = 144'hffecf0da09b40847f26ff93f0c1e0cb0ff2e;
mem[1084] = 144'hf94e0626004afbd50c40fa9708e109ad050e;
mem[1085] = 144'hf28a0068f192f984fd3ff9260c530dddfbdf;
mem[1086] = 144'h0bce0da3fa19060bfc2cf7d50ee50d78fe3c;
mem[1087] = 144'h05640b5804b0fb87f8bb077c04cdf0d40849;
mem[1088] = 144'hf1edf9220071f79102a00e34f97508ee0029;
mem[1089] = 144'h05e007050a5ffe63ff5ff83202a2fe83086a;
mem[1090] = 144'h0236f4e4f84bfde509bcf0d7ff8d0c70f991;
mem[1091] = 144'h0cacf0deff8d04a5f9e60f5e09e0f86af0fa;
mem[1092] = 144'hfe6d09c503e7f85bff48f553f5950737f050;
mem[1093] = 144'h0d6b04200a920b270021f990019cf42f0faa;
mem[1094] = 144'h05e2f82afb9fef5afbd40c2a073e0e09fb1c;
mem[1095] = 144'h04200cff07f20c09fdab01570e310d30f2b8;
mem[1096] = 144'h0bb80293f788fd9ff0a0f450fd8b0659f1fc;
mem[1097] = 144'hfe3502730cdffd9f0c81f9c50a460841041b;
mem[1098] = 144'hf44ef7330dcaf13df7ba0c85f6d5f4a20d7c;
mem[1099] = 144'h01250402f925050003c3fa37f41804d90bea;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule