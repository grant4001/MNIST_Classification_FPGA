`timescale 1ns/1ns

module wt_mem5 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'hfc0001d5ffe3face04250005029ef6f1f28f;
mem[1] = 144'h0967eb4aff7fecb30710007dfaa1eace032c;
mem[2] = 144'hf179fecaf89e0d52fce3ff21070ffca7ff1b;
mem[3] = 144'h084cef8c025f0a25f525f1f00663f7bf04ae;
mem[4] = 144'h0d74fa01f99af3c3f4020c3af1eafdc30bbb;
mem[5] = 144'h0231edd401de010ff645f930ee82fda50572;
mem[6] = 144'hffcf03400ce7fb6203aaf5db0319028f0552;
mem[7] = 144'hf73e02cfeebb03be0336f7cff932fa7cfacb;
mem[8] = 144'h0168f17f0603f6ec02430a0a03e4039c0d98;
mem[9] = 144'hf717fb950815f793022aff5df8ceede907c8;
mem[10] = 144'h00d0f992ef01f361f940f0d70a3a07b80364;
mem[11] = 144'hf0f4f1a7ffedfc5607740bd2f0a4f720fbb3;
mem[12] = 144'h01a2f376f9c5f345066d03d3fb2d0a58f829;
mem[13] = 144'hf46c02d8f9b9eeea045af978065202f6078f;
mem[14] = 144'hef41ff8b01e104710aaaf22207950ad9f4cf;
mem[15] = 144'h092ffcebf0fceffd04bcf705ee8df6c7f339;
mem[16] = 144'h003ffd86f8e5f8e8fcd3fbdc07b709e00cdb;
mem[17] = 144'heeddf31df360eb9507b303c4fe1e08fb0787;
mem[18] = 144'hf9100aec041efd14060efccb04fdef93fc9a;
mem[19] = 144'hfd4002760339f09ffa65f77ffe0d0725fa5a;
mem[20] = 144'hffe6f5d1fb2a039200e4f1ddf93a097dfc15;
mem[21] = 144'hfafffe30f8b908ee0496f42fecf1f25ff79f;
mem[22] = 144'hf4fb0cc0f3aaf4f2fbc0fb5cf930f742fa4a;
mem[23] = 144'hff3effc8f3a20b3bf6adfbaceeaa0744f98d;
mem[24] = 144'hfb31063ffeda048e0db30cf8ff930c7bf20f;
mem[25] = 144'hfb2af1b40996ee2001760a5cee59f60f0d2f;
mem[26] = 144'h01b90b140a210bb70079ef0d0999011e0a76;
mem[27] = 144'hf88404ddeeee0156f0dffa8a0830084604cd;
mem[28] = 144'h06270d36f7c8fb3a01b00344fcec0a6d01a3;
mem[29] = 144'hf1ca02c9f71ff836f0a40a4bf5acf786fca8;
mem[30] = 144'hff6ffbe6019a0481f0bf06f30cb4eff6037c;
mem[31] = 144'hfba6f61ffe1aec8406ca094e05d2f379ed09;
mem[32] = 144'h02be0db2f7dd0bc8f51cfb3aff3bf20bfbd7;
mem[33] = 144'h099204ee0bdeee46fae8fa4d0270f968fbb7;
mem[34] = 144'hf49807a4027d05e6fe8509d40500fb9c0309;
mem[35] = 144'hfd92fff7fa1f02d4f986ec7afedcf330ffc7;
mem[36] = 144'h086c01e5efc705edfc2dfe9cf68cf094f75b;
mem[37] = 144'h0014fec8084ff4ea07b8f46af1760814fd50;
mem[38] = 144'h069a04ce09c3fc91ffdc0248041302fa0982;
mem[39] = 144'hf331033afbccf321fd8dfcc10708077cf288;
mem[40] = 144'h011b0caa0d18f60d0ae8f458f88c0811ff33;
mem[41] = 144'h05b3f9d90576fad6f7f0fb7907700d57f18b;
mem[42] = 144'h0368fbdaf65c094c0b64075bf86504caf7fd;
mem[43] = 144'hf07eff1f07acf777002d071ff48cf537068c;
mem[44] = 144'hfc120517fbc509400d17f4a8fa69fee3f88d;
mem[45] = 144'h04a00199052ffa190b4900edf4d0038cfcbf;
mem[46] = 144'hf13e0746fd4700f5f6500a32005401e7044d;
mem[47] = 144'h08170494f80a057f0cf107aefd49fe64f642;
mem[48] = 144'hf2f50a160c2df43701ad0171f8b3009cef53;
mem[49] = 144'h0380f7990ae00c56ff89fbba0184ed71f768;
mem[50] = 144'hef11fad9f0760d8dfea10541047f06cf0479;
mem[51] = 144'hf6220dd7097c05d304700b3cf310f2220d1f;
mem[52] = 144'hf258f1bcf5dc0485f54e0492fb0ef6050679;
mem[53] = 144'h03adf1b50110f04bfc85028af7cc069200bd;
mem[54] = 144'hfca4f43d08c704a2f68c0a4f0c440300fb79;
mem[55] = 144'h03f60b8b0592edc7edab0c7d066b0691f380;
mem[56] = 144'h0790f9edff66f8a8fcd8faf5f70a06420b2f;
mem[57] = 144'hf1de09030d34facf0376f1af0a190d7102b5;
mem[58] = 144'h0d37069ff0dfffb7f020fcd1036e0193fe39;
mem[59] = 144'h091c0f3a0e2805ba0ebd00770de7f3d4f1a0;
mem[60] = 144'hfd3d0bb1f1abf7d703defeca01780d07f280;
mem[61] = 144'hfccbf283fe5a0918eda5f6faf86e07f8003b;
mem[62] = 144'hf6dffa8c02e1090cf703f89af083f2e10cc0;
mem[63] = 144'hfc4d0bb9f1b1f44802d70334eda4f00ff89a;
mem[64] = 144'h0aaf01b8fe3c05e402f8f847fb88f26000a2;
mem[65] = 144'hf289ee59f34d0117fd2bf3770344086b064f;
mem[66] = 144'hf3e0060102530fabf3eb0519fc43fcfe01a1;
mem[67] = 144'h0744fb740b0308ed058a0a0208e6084f0209;
mem[68] = 144'hf3cf06e20f2304c705d7f9c503a0fdc9fa8a;
mem[69] = 144'h0f680543f46e0da0f2b50e4fff7feff9f193;
mem[70] = 144'hf226fc6e05d00195fd1fff4b0615f0a002dc;
mem[71] = 144'hf6b50d98f9ba0e1809c9fae3085d0a680f96;
mem[72] = 144'hfa1608ba062c0932f6b1073a032af71406df;
mem[73] = 144'h07bdfb5bf5c1f79ff2990c5e05830836f714;
mem[74] = 144'h07f80a9009cff5f8f8a0f09cf91303bcf11c;
mem[75] = 144'hfdb1f1530e8002a3fb70f335fc9a007a0b07;
mem[76] = 144'hf868fec2003afb82fd63ff54f029f9e9f90e;
mem[77] = 144'h0190f4affd5008330f170d3707fffc0f0665;
mem[78] = 144'hfb22ff29f552091e0e2b004908aaf55df83c;
mem[79] = 144'hff5c00a40194f6a80166fc650c25f338fbf3;
mem[80] = 144'hfb4bfb51083ef7d1f4980f10fa31009af7c8;
mem[81] = 144'hf04f0054f314fad50bfafc30f481f3d8f877;
mem[82] = 144'h045cfc95feecfc7bf74c0763f71c0d37fd5c;
mem[83] = 144'hfd4af8ffff06013af08d010904210de4f234;
mem[84] = 144'hfdcafb8ff919039c0541f0d80db00e6706ed;
mem[85] = 144'hf059fee0f52608f2f0edf4dff313000cf2eb;
mem[86] = 144'h0aa2fe25fe8f0358051502bd0ada0be6f181;
mem[87] = 144'hfc1105820e710761f59bf6aaf46e0874fa31;
mem[88] = 144'hf65a0c59fc78fa1bfe25083f065700500774;
mem[89] = 144'h0dbbf517fdbffb13f7bc0a57f6ad022af544;
mem[90] = 144'hf82df8c6ff1d01840218fb58019bf69609d0;
mem[91] = 144'hf8fd0c67fb3f087cf9a8059f02b9f287f397;
mem[92] = 144'hfbe5f13bf284f0f4f505f1050b47f0f30f42;
mem[93] = 144'hf214f35f0c5cf8c3f6570bab04050376f96f;
mem[94] = 144'hffd70c7b08ad0ff9081ff33d06af0b19f065;
mem[95] = 144'h0d58faf0f49af45a0292074efb0fffbe063a;
mem[96] = 144'hfd11f4270cd0f1e9f1bd06ecf7010665fa76;
mem[97] = 144'hfe190eb8f01001e2fb18f2b600220dddf778;
mem[98] = 144'hef23eb2efbcffd07e37aecc1e2d4f9f4f363;
mem[99] = 144'hf29dffd0fb92f237f6bafeaef1900890f4d0;
mem[100] = 144'hf358003affcc0b27fea802d70b8ef0b7ef58;
mem[101] = 144'hea75efaae71ef770f67ff71de602e0230439;
mem[102] = 144'hf23101b5f11d060bf887f525f91c0b3deee9;
mem[103] = 144'h008e0b6cfeeaf852ee9902aeee08f8a5f488;
mem[104] = 144'hfa17049cfd46f901034bf1860267f419f9c1;
mem[105] = 144'h0df4f9d20c4cfd690573fc34f27defe7fd47;
mem[106] = 144'h000eeb9f005307e9fa32fdff0a4607400549;
mem[107] = 144'h08c30e49f7cf00f2fd62fd8307fef6760981;
mem[108] = 144'h004ef64ff3f9e999f7fef4ef03ef0804efab;
mem[109] = 144'h0a5e0881ff1b0346f31c0878095cf59a06f5;
mem[110] = 144'he47fe237e6c8039d055206990103f1f4feeb;
mem[111] = 144'hfd98f9200d1307c30cbff4c900bff13df52d;
mem[112] = 144'hf68afb4af18bf64af250e7f6e90efac4e973;
mem[113] = 144'hf338fb2c02350d460271f6f9eb9a0538f4a1;
mem[114] = 144'hfe3bfe9c07f7058efd15ee80ec3609120145;
mem[115] = 144'h0226fbfcf21e0bdf0c55f8b6034dfd65001f;
mem[116] = 144'hf1f6facff01007c1fb86078e0f13efaff647;
mem[117] = 144'hef63e98af600ffa3f0aa002df175f1abfcbd;
mem[118] = 144'hf2c00d1b0deeee720d16f8a6fef8f8320092;
mem[119] = 144'h04710588f34cf3ef0d1b031400950740087b;
mem[120] = 144'h07fef390f6f7fbf5f727087206eaf25d051a;
mem[121] = 144'hefc1efeb04a4f2910870f083026207e4f947;
mem[122] = 144'h027afce400faf89b0882fdfa027ff969fe72;
mem[123] = 144'hf360fb500e3405b5fdd2fb680ed1fdcb05e5;
mem[124] = 144'h0849ed91f789ea4507af0825070e00e3e663;
mem[125] = 144'hfd5dff4cff9d0e8301d4fddd08850e5ff773;
mem[126] = 144'hfeec03d5f6d9fcf3ee2c03520a6b067af788;
mem[127] = 144'h0de209130b75f0c2f633fdeff7c9f577f72d;
mem[128] = 144'hf111f8f3f0f7ed2ff05ff863fcc2f70ef8a3;
mem[129] = 144'hfe9df528f5e206340885f182012007620c60;
mem[130] = 144'hf663ff1cfe6d0194ea63f0300483fee0f37f;
mem[131] = 144'hef770cfaf54af6f406d900e4001afa94009a;
mem[132] = 144'hff4b0bd1f3a80510f89dee40f5b40113f871;
mem[133] = 144'hf296d91fed58f1e80295edb7f214e85401bd;
mem[134] = 144'hfbecf03defda0e2c009e0bf805c704e2f9dc;
mem[135] = 144'hf77a00a50b2a0e48fa230b200314f416efe5;
mem[136] = 144'h0ad8ef6806dafb49f186f18b03ddfe9ff286;
mem[137] = 144'h0842f85404b3feb00479f977f082fcf40636;
mem[138] = 144'hfc720c2afe21fc78ebe3faf4f0b20e82f5c3;
mem[139] = 144'hf58002910b1500d2fa62f3ecf5050b00f40e;
mem[140] = 144'hf5d7f866f63c003df96902dc1212071bfbef;
mem[141] = 144'h06befc39f42a00d8f03a0b5df734f80c0b1c;
mem[142] = 144'hf38bf36afeca0d2904a1ea46f3c0ee4ef753;
mem[143] = 144'hfa420f36f92a056cf58f0514feb208c4f335;
mem[144] = 144'hf2a3fff7fe1cee57eec2f754e591e51bee5f;
mem[145] = 144'hf25305e8f0e0027beedbf16b0009ee5b075e;
mem[146] = 144'hf946f185069309bd0203fbe3e73f0cbff771;
mem[147] = 144'h0dbdfb5b0561fe980097f0370d79f40f0025;
mem[148] = 144'hf4e4fdcafb28fcb70994f5fa0d28f6b00aa0;
mem[149] = 144'heac5f8570874ef6a0720faa6fcf0e961fa40;
mem[150] = 144'hf55ef9d4075ef2110d54f272fb6f0299f4a6;
mem[151] = 144'h0456f26df1a50a96f34902a1074b0ae0092a;
mem[152] = 144'h0e50f4f708c804d0fb12f09c0e7a0ec30e4c;
mem[153] = 144'h0491f5f6f3df0ab8f070fb27f1effd440916;
mem[154] = 144'h05d705a6034a0c04f45efdebf419f4bef966;
mem[155] = 144'hf796f07afd2bf265f78afe8009c00ed504c3;
mem[156] = 144'hfae1ed0aed1ced74f9e80aa7fb32033aef91;
mem[157] = 144'hf31ff980096ff0760d96ff5c00580b42f3fe;
mem[158] = 144'hf79409e1f66dfb88f0e9ef1c009d0d93f948;
mem[159] = 144'hf028fb5ef855fcbdfae208ed0c130ceffbe8;
mem[160] = 144'hef00f1ba0beb0cf5f0a507f0f488f6e00e2e;
mem[161] = 144'h03e90ca5f2de095ffbc5f8d9f3750599f4af;
mem[162] = 144'hfbe5fe660dad023eff4401a209f503d6f437;
mem[163] = 144'h05d4f37802aef9aaf21a0765eff60199f394;
mem[164] = 144'h0703f37c08bd0f67f7ea0e36f32b07d500ae;
mem[165] = 144'hf45af344f61afba403fd0055fbe304cdf847;
mem[166] = 144'hf894f53902360b390bf10b1a06de0926032e;
mem[167] = 144'hf5b60785f99d03f008b9003d047801890b0e;
mem[168] = 144'hf73703bafdd7fc9df3db0cacffdcf3d1ff06;
mem[169] = 144'hff4ffb7ffb5504d5f23b03830c060c640356;
mem[170] = 144'h0cb0fe9af47f09dcef8206cff4e300f10073;
mem[171] = 144'h099df706041c07b10b60fa2705f6fc80f134;
mem[172] = 144'hefc6f029ef9604000a5901b3ee530a5708df;
mem[173] = 144'h06bb06690b9f05f7ff51ef490eb00d570491;
mem[174] = 144'hf751efe6f5980bbf0decfbc5f818fa86f56d;
mem[175] = 144'h0d61f459fa7efdb4fdecf65d00730df002c6;
mem[176] = 144'hfe02f7ac0352f2d20575fcefef5d0c6b09e6;
mem[177] = 144'hf8b705f20948fac9f79af43f0620f446ff60;
mem[178] = 144'hfd35f9b00a0ef47ce399fefefc1805baf9f1;
mem[179] = 144'hf72ef78704dc0709f3c60a520573f614f4d4;
mem[180] = 144'hef6a0a49f9c002b4f6eff2820a0305bdf30e;
mem[181] = 144'hfe4f0593f53b0afd0216005ef4b9fb77f60f;
mem[182] = 144'hfe23fa6a0cdef511f08f092ffbb108b40023;
mem[183] = 144'h00ca0178f692f69106af004bfd6cfb05f28c;
mem[184] = 144'h08f80943f207ffebfd770581f3f10e0302b9;
mem[185] = 144'hf6c4f626ee750c3d0d0fff53f6a1f5cbf661;
mem[186] = 144'h0ab9fe0408110ae6fe2902000858f1f1f7ad;
mem[187] = 144'hf39005e4f0f706e10928f2ec0a800ab3f8cd;
mem[188] = 144'h0496f2c9f5abfb02f219fdb3fad5e4e80727;
mem[189] = 144'hf6f1f4ea0993f50afcaff5f80858fe3df107;
mem[190] = 144'hfbdbfc4a0d8ff7b0f376fc7207f3ecc90b3d;
mem[191] = 144'hfabb06fe07cc09100b86fe7a0c0904cf06a0;
mem[192] = 144'hf0b9f82bf85506c2fbceec390801efa9f511;
mem[193] = 144'hfffc0b190d86fff30203fcc30c27fa4ff37c;
mem[194] = 144'h08940b4cf143f78a05ebf3eb09c8f00ffb12;
mem[195] = 144'h0818f4edfe6509a7f0550ab9fcbbf3c0fd0f;
mem[196] = 144'hf59bf12301b5fb4b01f10ea3f381fd02f474;
mem[197] = 144'h08f0084b0209f4f5fa74f8e1004afca2f2a7;
mem[198] = 144'h0aecfb89fcbf09d30545f3cc0c2ff8d90b23;
mem[199] = 144'hff1cfb3d0bb80cd10879f92ffdfbfaf6f58c;
mem[200] = 144'h0822fe5805410dacf2f2f2f9fd2f09810333;
mem[201] = 144'hf97aff33f7cafe410a89f61ff258f4daf008;
mem[202] = 144'h064ff925f4a20e46f1a70fadf87c0257f80c;
mem[203] = 144'h0bf60d7efd6b089b0d6f00110f9af1b0fb45;
mem[204] = 144'hf9c1050f05540309f6a809f2f3b0f0390b92;
mem[205] = 144'hff69f10109b9f3a3fe170d93f2b20d7b0f9f;
mem[206] = 144'h0f71f7060817f92cfbae0434f7af0061f05e;
mem[207] = 144'h0fcff75cf4c10d29f1170e14f44804cc0613;
mem[208] = 144'h0487f185f1fa05790d15ff57ffe4fddbf423;
mem[209] = 144'hf22af8adf78904e5f2e8f671f70ef920009e;
mem[210] = 144'h0d8fefcf0ec5fc7df0400531fda300de0d6b;
mem[211] = 144'h04e009f5092d09110ecff0e505c108510608;
mem[212] = 144'h0b21f721fc23f57c03b2fb050c78f785fcee;
mem[213] = 144'hf42602880790f95501480c5af393fe650370;
mem[214] = 144'h09e20885005402bdf268f49ef81bf2c0fcb0;
mem[215] = 144'hfa2d03320baaf7a60bc3fe910ce5f0b1f011;
mem[216] = 144'hfaba0945fd92fd6b06850290fccf0ec2fc2c;
mem[217] = 144'h0d010dcf0adcf5ce0ac502fbf923f01b0a80;
mem[218] = 144'h06f8f4c00373f8a5f9e90eacf208052a075a;
mem[219] = 144'hf97701befdc20a3af730f12a0460f9a1f065;
mem[220] = 144'hf0cdf5a2fe30f2e4094dfb920169f040f829;
mem[221] = 144'hf51cf358f35ef10a0c46f6e600eef36c0062;
mem[222] = 144'h02c7f83cfe70fd3c005ef8700b500a27f4c5;
mem[223] = 144'hf729f14b06bb0f080fd80bc6066f09420e81;
mem[224] = 144'h01520aadfed10ce50229f2ccfc6d056c0bf2;
mem[225] = 144'hefeafeba05bb0899f18cf7f809bd07ccfbfe;
mem[226] = 144'hf430f6730c69f0bf00f7053afb16fd0e0c6a;
mem[227] = 144'hf9100424fe950c090a970d21f255fea008fc;
mem[228] = 144'h0a8df45c07fcfa44fe610c1e041c00b2f50a;
mem[229] = 144'h0c72fb1e0c380ea0091ef720f73103480d8e;
mem[230] = 144'hf1890137093df8c60f3007ea06c30363f1a5;
mem[231] = 144'h0766fedf0b7d0b3505dd0338fa65fa27f91e;
mem[232] = 144'hff5df0eb0db4fd63fbc2fbfff43a0d51f2b8;
mem[233] = 144'h0f04faa90ccafd15f77afa340519f74e0575;
mem[234] = 144'h06cc04d2fa42f189fe96fe7d0aa3f44cf846;
mem[235] = 144'h04020ad5f3f20c82fd8d0a7a0eba0b63fca5;
mem[236] = 144'h0babf470043f07d8f5550b3df028fac60eac;
mem[237] = 144'h086d0a00fcc402e3f3b9f8050d39f595f1be;
mem[238] = 144'hfc3f0a12f9ab09740bc50354f46c06bef3cb;
mem[239] = 144'hf98c0997f274015dfd100e17f7e705fff1ed;
mem[240] = 144'hff54fd45fd92f6adfd3b0518f6baf0710021;
mem[241] = 144'h08280dfef751f93f072aefd60a270e65f9c6;
mem[242] = 144'hf80c0c120464f87c0f8f0d34081f0404093c;
mem[243] = 144'h011e05170c9cf2b5fe28f30008350733045c;
mem[244] = 144'hf676f9a20f83f8180b94f8d5033809580e37;
mem[245] = 144'hf1510cd0fb740ecbf4c8081cf55cf37e0145;
mem[246] = 144'hf474069cfc9f049c075ef554f3bbf4f40feb;
mem[247] = 144'h051303e3f77cfd3a046c07c500f4f977f028;
mem[248] = 144'h0eb6f0fd07d7fff6083b089ef99600d7f857;
mem[249] = 144'h0f16fcaffa67f36c0f950b9d03f80991f090;
mem[250] = 144'h04ecfff6061ff4f80bc0f226f3e40081f053;
mem[251] = 144'h09e50d77fc8ef1c10d7d0067fd690b48f4a9;
mem[252] = 144'hf3810552fad40c2afe38f909f67eefccf91e;
mem[253] = 144'hf7cbf40a07ce0e90025602bcfce708a30804;
mem[254] = 144'h04a6f3020a750081f10a0a510783f6ccf5aa;
mem[255] = 144'h0a810a660b540da009ef0252f5cb068bfebc;
mem[256] = 144'h0051f0aef34200dafbe7074ef18307e4050d;
mem[257] = 144'h051e00f8f7ddf375f74809a607bd01dcff59;
mem[258] = 144'hfba8f6cbf0490c13fa220a1ef8af0097f224;
mem[259] = 144'hf1c60531f22504740f740adaf0fff32a024e;
mem[260] = 144'hff8df81cfe4e0c870cba04c4fd47085af426;
mem[261] = 144'hf6e7fc1cf6ab08f4ff7ff7230378f51802c3;
mem[262] = 144'hf594febaf4d80b40f62802a8f9a0efe7f05e;
mem[263] = 144'hff2f02d2fb44f0cbfc30f9fb006c07390827;
mem[264] = 144'hf243fbfdfb780bb8fec10a19051f0e99f84f;
mem[265] = 144'h0444fbd9f2bdf31cfa65060ef030efb9fa2e;
mem[266] = 144'hf8ea0d62033df264043b0b56099401bafe5a;
mem[267] = 144'hfc43f7ae0206f0cbf0f0f5e6078a0218f4a4;
mem[268] = 144'h0a20fd3705de0570055f014dfb4d01c8f3e0;
mem[269] = 144'hfac8046e0843f2e5f7e5f979ef0eeeb8f05f;
mem[270] = 144'h0aabed9bfe53fca0ffe809af0b130e9508f4;
mem[271] = 144'h0efafecc02dffcc50e5b0c6bf861fed5f19d;
mem[272] = 144'hf653f073f960f41f0a0ef8980943f8fb0116;
mem[273] = 144'hf096004e00a9f40cf553f18006c9f67f0edf;
mem[274] = 144'hf42ff2df0ed8ed5dee82daf2f13ef3aafd10;
mem[275] = 144'h042e00ce03a1feb908a2ff5d025bfd450de4;
mem[276] = 144'hff7f070cf21c0bd80957f0d8ff81fa59f712;
mem[277] = 144'h0129ffd9fe0b0a2903b5e754edf60193082c;
mem[278] = 144'h09acfffe00fcf8d60021f966fd5cf86df2cc;
mem[279] = 144'h05f50a55ff560baefd1d0b41f7d10c370b31;
mem[280] = 144'h049ef8d0fba70d4c00930a70f275f703ff55;
mem[281] = 144'hf1c5f93302d0f31504390708fb0d0ad00735;
mem[282] = 144'hfec501d5facb0533f588f3350129f33ef569;
mem[283] = 144'h052ff0270142f2a8fe6903280e41f6180bf3;
mem[284] = 144'h0e6607f7ec43f5f20e44f72b07f20bfff6f7;
mem[285] = 144'hf3fa02baefe7f7b005fefc5f0c4aef400b2c;
mem[286] = 144'hf1c4f3080b0d0158f5e8fcbb021f050deefe;
mem[287] = 144'hff40019506daf438f10707630e4d054cf6c0;
mem[288] = 144'h000300abfde8efbb0450f93efece0203094b;
mem[289] = 144'h057bf9d2f5b90e3b031df15709f10ceef19c;
mem[290] = 144'hec1af85bfc52fa590393f7ec0008ff27fc93;
mem[291] = 144'h0d11f90109a7fa47fef5f02fff7b0176005a;
mem[292] = 144'hf4a303f1f3330e76048bf0e2ff58fcd2f0d2;
mem[293] = 144'he000ebeef97ff80ff311e714e48cfdfcfafd;
mem[294] = 144'hf68ef46a02290a96f8e207a9f9370b12fcb7;
mem[295] = 144'h0c19f147015a0922fe2ff3560df5f19a08ea;
mem[296] = 144'hfc5ef9d6f4dcfe8ff8c0fe7e0cbdffebf6b0;
mem[297] = 144'hf3f7010cf67b08b90a1dff090b86f9f6ff84;
mem[298] = 144'hfcec0be4f4cbee6ffd1f0ceaff1d0c270acf;
mem[299] = 144'h04af06e9f99a07a7fd97efddf4a701b607b2;
mem[300] = 144'h0031fcbef18feec80f2afb270446070aeff7;
mem[301] = 144'hf5fef94a0ae4ff2eef1bffb8fe2ff0990b3d;
mem[302] = 144'hfcf9f9df0abff09f060ff7e1ef53efa4f745;
mem[303] = 144'h0c43f927f3d4f10ffcd207490e7bf0f105d3;
mem[304] = 144'hf9f503aff61105e8ec44fefff429fd7a07af;
mem[305] = 144'hee00f416fc4e0120f408feb4ed3cfd6af561;
mem[306] = 144'h0a780971fc9b02e9f685f57008910b30fca4;
mem[307] = 144'hfea3f2c9f9cc023ef3a4f3b300960b2ff91d;
mem[308] = 144'h0d1d0f34fab50db9f33c0b5c05c50f900c74;
mem[309] = 144'h0a4cf842f6c20b51f68a0d30f8e1ef780c90;
mem[310] = 144'hfb1005290a330c9b03450797053bf5d8099a;
mem[311] = 144'hf729042dff230d1b016dfa13fec70d9df815;
mem[312] = 144'hfbe2f6c7052a047df454fd4b0ba2ff15fb10;
mem[313] = 144'h0d2eff72fe960cabfc1a000f0923f53df015;
mem[314] = 144'hf1430a3ff7d6090904140d0cf27803360431;
mem[315] = 144'h0313f0e4f7450a000ea0feeef3f30dfd0007;
mem[316] = 144'h0a26ec83f3cef27f0864f1be0b8208ee0ac4;
mem[317] = 144'hf00c07a8f434f7320e20f3730d47018dfad5;
mem[318] = 144'h0180032b0e30fe48046efd68fa9b012ef768;
mem[319] = 144'hf5c0016604cefa06f31bfc540ea70a3cf1c2;
mem[320] = 144'h055bf2ebf1f7fdfc0d810ab6076cfcdcf7ad;
mem[321] = 144'hfd28f415ff5c06c001fbffe00c3b006a0b47;
mem[322] = 144'hf6cb018000100c2e0726f51df667ef8a0ec7;
mem[323] = 144'hfb3f0a6200f2fac8f61102aa07080d0df607;
mem[324] = 144'hf8defa68f94f0bb2f23bfd5d01e50ca6070b;
mem[325] = 144'h0aac06a40adbf7e00bd0ee6e0978fce00c3b;
mem[326] = 144'hf90bf9e00f670c4dfea300d50971fcd5fc9f;
mem[327] = 144'hf4c403210a6c03860574fffa0ae70b0f03bc;
mem[328] = 144'h0f4f0c01f5a90862f6a10394f33fff91f632;
mem[329] = 144'hf6fb002f098cfddf013bf14df754f913f9c9;
mem[330] = 144'h0765fa8efe90f7a2f5c0fb95f2bb06eaf412;
mem[331] = 144'hfd8e0147fd63f5bb0661fa6b088e02830ddc;
mem[332] = 144'hfc78ef9f05a8f13e0144fae0eb40fa7ff0fc;
mem[333] = 144'hefe9060bfacaf677fdde06c0f37c060df8b3;
mem[334] = 144'hf789ffb10c2d06eef3eaf83a041302980944;
mem[335] = 144'h0ba90bf40a24ff2b095a0a84fa7eff37f8d9;
mem[336] = 144'hfbff01840e71096a0cdaf5b9f446fc8efb52;
mem[337] = 144'h04e9f72fefa60adff1e807c40d3efdac0f25;
mem[338] = 144'hf6fc0a0201a5fcabf593f039fde3f3f7f79b;
mem[339] = 144'h0d50fa100bb5f69b0a8c070bf8c2fb36f6e3;
mem[340] = 144'h0e6efd760d56f5300ad301fbf6860788f686;
mem[341] = 144'hfdf609b300fc0943f5b207daf3a10a81f931;
mem[342] = 144'hfd9c060afaef0c2509230bc40d3500190820;
mem[343] = 144'hf89cfdc4f6570f8e00b50e4effad01f4f1af;
mem[344] = 144'h0088ff950c3efb2c055a0d1805effa4f004d;
mem[345] = 144'hf706f606f0bffb4d0054fafefc90f33cfead;
mem[346] = 144'hf269082df7690d170f45f0eaff7608d40942;
mem[347] = 144'h0f53f1c701230aa50d41f60807040e300722;
mem[348] = 144'hf929f2ee0860f383f79c07baf1cbfa3607ee;
mem[349] = 144'hf319f28f0a41ffb0f2ca05fdf2f701a40d54;
mem[350] = 144'hfd08077ff4e70c9ef8e50c37f40ff71ef1cb;
mem[351] = 144'hf806fec7f239f884f0a7fd08f19b00f8fcb2;
mem[352] = 144'h0b6ef9480625fe19f88101a105e00d950041;
mem[353] = 144'h094c0597078d050c0ccf04540710fa4bff7f;
mem[354] = 144'h0cd3f1140e69febbff96f3c9012905a9f340;
mem[355] = 144'hee60029500a3f7a4f8dbf0a2f506fab4fd9d;
mem[356] = 144'h0467fe44ffabf3a4f8b90567f948f4d4f93c;
mem[357] = 144'hdd1aea75fc9dff95079dec49fdbd01990913;
mem[358] = 144'hf2a00baeed9cf506fd40f5980acff348f961;
mem[359] = 144'hf219f45cf2e0027ef7f503e50624f375068b;
mem[360] = 144'h0431efddefc4042bf7bd073efda9056f0530;
mem[361] = 144'h07d30a670d0106fdf6360382034ef484feea;
mem[362] = 144'hf34ffa9fef54f7130a8502bc0aaffc7c0137;
mem[363] = 144'h04190bfa0179f12f02e00002f68a0103f40a;
mem[364] = 144'he986028af29cff9d0e78f590078cf2d0e871;
mem[365] = 144'hfc4106f9f2f0f0df06860a85f65ffccbf0c6;
mem[366] = 144'he309fc90f79dff21092bf08ff5ccfdfb0a39;
mem[367] = 144'hfec80b82029f0155052ff3c2093601a70a5e;
mem[368] = 144'hd20adaadfc80f77de925f35ce7b2f7480831;
mem[369] = 144'hee95fcf10166eecbfb7ef1ecf128fd2905f9;
mem[370] = 144'h0640f4100b23ef98e4c9ea20ea76eca70952;
mem[371] = 144'h0be7fec408f5f23f06c6f4ce066df2bb0199;
mem[372] = 144'h03570cc9027f04410c620e2d02d9f17302e0;
mem[373] = 144'hf547fd78f607ef0a0182fffd00be0116059b;
mem[374] = 144'h0622047bf08fedc1f1b307c106710251f8b4;
mem[375] = 144'hf33102cef0cdfc36fb24f656fba70579fa56;
mem[376] = 144'hf39c0639f1b7f536f2c50b8b0aa4f884fe3f;
mem[377] = 144'hfd6d06e4fd10ff03093cf7b4eef0f95eff11;
mem[378] = 144'h08d20b60004e0d8df14d07dcf1f5f04bf36d;
mem[379] = 144'hefc9006e038ffe7107a5f64df6a4f56df554;
mem[380] = 144'h083f0569f7a8f801ead80358057a04d5eb94;
mem[381] = 144'hf1deefe80866074c000c090dfc33f8ca085e;
mem[382] = 144'heb6e02b10daafb750bedf8b9022d09d100fa;
mem[383] = 144'h0a0ef1e2f7c7fe59ff620d7ff33bfa180182;
mem[384] = 144'hf560027aece90a5ff2f4f45df03de909ed0f;
mem[385] = 144'hec5ff818fa49064d005a052af800f2710741;
mem[386] = 144'hf65def7dfebae856fa82fae4f15ee107f0b6;
mem[387] = 144'h027b04250188f381f318f6ac0a9f03770c7b;
mem[388] = 144'hff55016ff18108bf0168f176fe55f0c80250;
mem[389] = 144'h0341f7b8fbc700f4f22ff538f1140a70fa1a;
mem[390] = 144'hf285fe44fbd9ee10faeef1b80470edac0059;
mem[391] = 144'h0867eed10750f6a7f80003980bf0f09f044f;
mem[392] = 144'h036402e107edf86d04c8f42af5ebfe0a0da2;
mem[393] = 144'h0680089ffcaf01aefd07f37cfd6702160268;
mem[394] = 144'h09c3f1880afafa720b390cbf0477f70a0133;
mem[395] = 144'hf27c06810526fbd2fab5ef0001e90497f467;
mem[396] = 144'hfa6cf01afb0bfb0ef48f0935111202880043;
mem[397] = 144'hfe98f9b3010c00220a30fb61f23cfce4fa1c;
mem[398] = 144'h050a044d0c9506fdfbf4ecedfb59fd8fedae;
mem[399] = 144'h063e0647fc160961027dff63f3850318f96c;
mem[400] = 144'hedddf7b3fbed0bbcfb8f004ce965fcdbf155;
mem[401] = 144'h0483f77cfa8b057701aaf2ba031fec540237;
mem[402] = 144'hfa9ef1370bf801f6fc0df4d70610f7250e05;
mem[403] = 144'h09abf7c30b66f94606d80656f448f61cf985;
mem[404] = 144'h0845fd1af850f0e1efa3f1f5f1fbf7b3f1ec;
mem[405] = 144'hf57af4a7041b064ff4e3ebaa049afae10601;
mem[406] = 144'h0785f34c0e4c044a06c40112048a060d0c6d;
mem[407] = 144'hf46c059e09260853f6810445055eff27f9b8;
mem[408] = 144'hf2530d9ef140f67df5410bbd046b050c07d3;
mem[409] = 144'hf2cbfdde04f0f463f9fc0132f06601ac0136;
mem[410] = 144'hf55d016bfe3607fbf980fddbf2f1ef52f7a9;
mem[411] = 144'hf659f385ffa4fd580646f753f06efdcdf08b;
mem[412] = 144'h060afbcf0497fd43ea1c0a750e2de78b08e7;
mem[413] = 144'hfab408b8f367fbd6f641f302f2c7f62df5e4;
mem[414] = 144'h001eefc3f6b60367ef66ee48ffbaff340a25;
mem[415] = 144'hfde002d50ced06bff6fbfd110c7e00f203f1;
mem[416] = 144'hf9dcede3fb45fb92f704f29df8f4f401fdad;
mem[417] = 144'hf37e009901e000b0f6b00859ef3800b20017;
mem[418] = 144'he75f0419fc7905bde956e21bf2df0a7909a7;
mem[419] = 144'h0b07f907fe0e0301f196088cfb990bb4f8fc;
mem[420] = 144'hf65dfddc08f1f7c1f671f3670a14f48cf589;
mem[421] = 144'he13aed4ff4210e42f107ee9be889eab403c0;
mem[422] = 144'h0a150985f015f97af96ff997014bf935f46a;
mem[423] = 144'hf116056c04d90d57fcbaf0d80a06efa2f6ca;
mem[424] = 144'hf11e05280c06fd41fba0fcca010ef667f06a;
mem[425] = 144'hf1290180f9a2fcf108d6009bff8cf961067d;
mem[426] = 144'hf28cf3d9fefaf2f9f6bc01f7051a01840db9;
mem[427] = 144'h0d21f82ff8b9f305f5e00b65ff76f34d0dad;
mem[428] = 144'hf4a109cff453f8a6f6550cab0125077efd7e;
mem[429] = 144'hf7330dab019902a80cf10331f4e600daf21b;
mem[430] = 144'hff7d08c3f6080da1f655f114f54403b1fe3c;
mem[431] = 144'hf1a70a9e0108f6420a9df340faf70437f001;
mem[432] = 144'h0130f14709280fac044102c1ea5f00930293;
mem[433] = 144'hf36ef8c605330a89f9cef244014cf722fbe6;
mem[434] = 144'h085e032ff186f97d0f35fc6001d2037f0eac;
mem[435] = 144'hf37e0600f2f5f4e506b702aef30cfc7703c9;
mem[436] = 144'hf3b20e6e0134f051f48f097f0ab8fba6f58a;
mem[437] = 144'h0eab0b5df252f216f414f8a605a1f1e50bd3;
mem[438] = 144'hefbcff8afb9df6aef4db0464054ef586f3a6;
mem[439] = 144'hf5b8f1cb061e0e81f2f9f2d6f747f3b7052c;
mem[440] = 144'h0171f8ec0898f90c013d043eff6a01250cd6;
mem[441] = 144'hf4fdfec0fcabfbdafb45f2b8fc08f2170f07;
mem[442] = 144'hf239f2e7fc580541f0b3f6e8fe56f9b1fbc6;
mem[443] = 144'h067bf7dafb8affb60e75f852f7370ce0f2f1;
mem[444] = 144'h09fcf1fef2b2f610f983f232f78cf5200f03;
mem[445] = 144'hf73404ba02f20b8ef85a0c590ed2f44cf30b;
mem[446] = 144'h0377f7210407fb98fec6f69dfa6bf97d00b0;
mem[447] = 144'hfaae09480dfd064bff58f843fe12f85af098;
mem[448] = 144'h0bba0439ff20fc32fde0f27dfb83fc4706a8;
mem[449] = 144'hfbe4f4b703370670f422051a03600304039a;
mem[450] = 144'h08a20916f9c00212f6bcf4770a75f0550859;
mem[451] = 144'h06690f1e0daff1f4f3ae0bce0dc5fe7af6f5;
mem[452] = 144'hfb4d02a60e12f76cfd23f515fa5905c90b66;
mem[453] = 144'hf86706540307f6ab06b4f24203900d7d0137;
mem[454] = 144'h09eff7e0f543f35a04e20093f8fdf865fe84;
mem[455] = 144'h0ce303a4f13ef51ff3daff6b0d2bf2b5efe1;
mem[456] = 144'hf52608c9f310fe61f2f9f362f976fc250069;
mem[457] = 144'hf63a076c0927f327f1df05890f36ffe60d0b;
mem[458] = 144'hf61ffdb70f2af8740322ff82fff2fdb8f0bd;
mem[459] = 144'hfac00924f997fe5b06dd0667f2f508e20e81;
mem[460] = 144'hf0d9f9860108f1b3f5350451008b03610d40;
mem[461] = 144'h0a6afeca0eabf0d80ed507e6033a0931f2af;
mem[462] = 144'hfd9506b0f4e40af00a1f0a1d0b800d800717;
mem[463] = 144'hf415f762086ff54501a5fa42f0800fb6fbf6;
mem[464] = 144'hfe7902defb770baa01760142fffd0bce041d;
mem[465] = 144'hf0140edeff0b0ee800cff837f94004aa0a17;
mem[466] = 144'he7f5f469fa03f929f18bff1dfda8f96e032f;
mem[467] = 144'hff96f850fcd1efbb0d27fdf806def530f539;
mem[468] = 144'hf152fafd00c3f7890a86ffdaf3fdf2400174;
mem[469] = 144'he257f815f6e906daf6e1f8b6fb5ef107033d;
mem[470] = 144'hf7bcf44f0a1ffab4f590fa24fdf903e10dfb;
mem[471] = 144'hf73907300ce5f4fa09b50182eff5f28d076e;
mem[472] = 144'h0889f13cfdf507c900eb09f10d9908eb03bc;
mem[473] = 144'hff1df5c4045c0d2ff62ef7e903350034fa82;
mem[474] = 144'hf7eb034df0b1094a0bd102c90a66fea40cc2;
mem[475] = 144'hf76b0b8fff5c06e5fc6606d40cb8006eef20;
mem[476] = 144'hfccc04faf1acf019dd7e08501b58e862e894;
mem[477] = 144'hef4c0579fc3508f0f1590a28f9a50accfb40;
mem[478] = 144'hf0940426f9f10095f98dfe4202c70664f22a;
mem[479] = 144'hf15d050f05680ff1fb350ec70902f3e60abc;
mem[480] = 144'hf86cf6dc01a6f4acf3a1dadbf010f419fd2f;
mem[481] = 144'hef18fc8708c70294f486eda8eeacf37508a0;
mem[482] = 144'hddc30450fe56fe14f8b2d9a0f95cf28b0f73;
mem[483] = 144'hff1c0a5a0000086301bd0d45064cf16ceff2;
mem[484] = 144'hf8a4ff6cfbf10ccbf22e04c80a590a71f531;
mem[485] = 144'he6c5ea9305ac033ff3e2f230025bfbafed3a;
mem[486] = 144'hf13a0b22019af83af8c8edd70ae5fc8a0701;
mem[487] = 144'hfd98fc3102080d4c0061f050070cf8b2068f;
mem[488] = 144'hf35af83101baf732fffb0c51f1c1f4c5068d;
mem[489] = 144'hf4b8f001049607d001760cb501320677f7ab;
mem[490] = 144'hec79fbb207c20bc102eaf9f2ed130b04f4d3;
mem[491] = 144'h07f6fd62f4eafd8107e7f9b900a206d902b2;
mem[492] = 144'hf50d087afa8dedecf326ff7a09430691e6bf;
mem[493] = 144'h0c37f7020313f81af2a40e0308b7f136efc9;
mem[494] = 144'hfe76ebe0ff590b9105beeeacf629fd8ef099;
mem[495] = 144'h061606240d9ef9e0f9ac0e8c04e6f3bd01be;
mem[496] = 144'he388f7690735f985f9ebfe96ff4ae8d4f0ad;
mem[497] = 144'hf343012dfaf10812fd3c05d5f42a0bc2037d;
mem[498] = 144'hfa1207abff84fb6dfee10555fa90f86501e5;
mem[499] = 144'hf9f20cc7061705c8f87ff842094108ff007f;
mem[500] = 144'h0f450f910ed9fbbf0db10fa0fa26fef3059d;
mem[501] = 144'hf78dfc4afa0c01e2fc78f0f6f0fa0c5c07b5;
mem[502] = 144'hfd0f08740c360341fc56f6af06380c70f4b3;
mem[503] = 144'h0f20f4bdf4530403f2d803a1f4950951019c;
mem[504] = 144'h08e9fa7b034df21a0392f4d6faba0536f0af;
mem[505] = 144'h0f150bfc0240f2e1f31008c008350dc0f8ac;
mem[506] = 144'h086ffa22fc12f0af03ee027b0b3bf369fd61;
mem[507] = 144'hfa4f030ef29d0600f476072ff3650d640ec1;
mem[508] = 144'hf05ffc10f43ff608f62707a4f10408f3f074;
mem[509] = 144'hf2ec0783f6f601e204baf7120b95fea9f6e3;
mem[510] = 144'h0bc8f9f8f61aff54f6b005ccfaeaf223fae8;
mem[511] = 144'h08a4f324fa24ff04f71ef072f06eff3bf04d;
mem[512] = 144'hf4270ac9ff85fd1a09d10a2ef98d047df436;
mem[513] = 144'h02def364fc4905d90e9bf278f16efdf5f619;
mem[514] = 144'h0420087e064c036a06cd066ef9b5ee37ff2f;
mem[515] = 144'hf39309b4f10ff331fd25049e00af08d8efe9;
mem[516] = 144'h028008a40307ef840c1b0127f71800bff270;
mem[517] = 144'hf44a06dd0188f2b106acee39fe220931f28f;
mem[518] = 144'hf207074b06e1ee94f391f6f205d6f7b107ed;
mem[519] = 144'hff0f0b4e071effdc02a4f783f0d80d920eb0;
mem[520] = 144'hfbf5f5d0f66df1cdf433f316ff3ef99804fe;
mem[521] = 144'hefebf66d02c3f92c001eff3907b5ee1006db;
mem[522] = 144'hf79a0c0701c2038ff5b4f3d1facf04fcfaa9;
mem[523] = 144'h06c5fd5a0861007ef25efdbb04790385049b;
mem[524] = 144'heb6ff92a0976f7c1033eeb1cfe02054dff8a;
mem[525] = 144'h0de8f705014107b50ab40e4c09cd04dc09fc;
mem[526] = 144'h0641f6fe08b7faf106fcf3d90a12013a0e20;
mem[527] = 144'h0359f6930bfcfda802c4f003fdf60df208b8;
mem[528] = 144'h0441f235f0ed0560ef5103afed80ffa60b76;
mem[529] = 144'h062c036e0c6f0ddbedbffbb2f47ef071fd19;
mem[530] = 144'h0376fd39fbb70128f0e2ef5df50909caf80d;
mem[531] = 144'hfa2a07fffae106640d6a029cfb41feaf01b0;
mem[532] = 144'h020af2b80e18048bf7ccf8e00b4df28cf014;
mem[533] = 144'hf921f50afcfd0dbb013afa1dfb5803e7fe7b;
mem[534] = 144'hf057f300ff24f2030db7f1830011ffd90606;
mem[535] = 144'h01280dc3038003c2fe13efcd096afa2dfbc6;
mem[536] = 144'hf9cc02a2f4e1f7aaf87907100fa3fa9c084f;
mem[537] = 144'h078809c7f641f82cf39cfc070c35f48efc17;
mem[538] = 144'hf8e4050e017306a400d0f1c9f2e2f4cffff2;
mem[539] = 144'h0406fefeffbaf198f6100959f719ff900de7;
mem[540] = 144'hf5a4ecdcf833047a0292f4ff07d203330583;
mem[541] = 144'h00d1fa4af4fff49bf655f3b4f7240c9c0e8f;
mem[542] = 144'h0c92ef2ef71ff1ccf344026c0609f1b00bde;
mem[543] = 144'hfc84fca9f8b0fa9e0627006cf44ef4420c07;
mem[544] = 144'h078a05bdfff600fa0211f9b9089f00f5f1d4;
mem[545] = 144'hf39f02380c09f1bffd03012503770c10f523;
mem[546] = 144'h0ee5f5d90e0f0d9af40df435ff7f0827f61b;
mem[547] = 144'h0554f82e0949f4d9002cf8c3f4f00b2801a5;
mem[548] = 144'hfe5bfc1c085a09cff11801990997f46f01f9;
mem[549] = 144'hf444ef1ff76f0f22f442064df89a0ce30027;
mem[550] = 144'h07dffa7df21401390e44facd0e22f953f9a9;
mem[551] = 144'hf687fc23026c0f160ac3fd6000ae0cb00b2f;
mem[552] = 144'hfc3a01c2002609bf090b0115f4ccff89f403;
mem[553] = 144'h06a3fd920cc1fee3075e0946f9590cc20b26;
mem[554] = 144'hf87bf79200f4fd5bfe94027804d9f860f0c2;
mem[555] = 144'h0099f4b001b9fec8fe4805930fc3f46affaa;
mem[556] = 144'h03efee6ffd5ef9e80828eeff04bd079af922;
mem[557] = 144'h0d8df8380e5e097a012b0ca10278f475fd60;
mem[558] = 144'h0a460aa60d25f3d6ff45026b0b79fdfcf1f8;
mem[559] = 144'hfbe90c68fe75f8ec0719f93af57ff24a0832;
mem[560] = 144'h0e080822f57bfa5706f9fa7802d504100ad4;
mem[561] = 144'hfbb8033201680f260716fd01f95d0ebcffa6;
mem[562] = 144'hf4c1f9aff894f66c0b2cf032f25e06fbffc4;
mem[563] = 144'h00c20e4cf034f3d6f207f8ed0c590405f25a;
mem[564] = 144'hfe41089cf38af2aefeed014df862f0fffb66;
mem[565] = 144'h07c4f254fec2f9b5f2c70a64f3ca0535f983;
mem[566] = 144'h0b84facc00720efaf066fbe4f0e70e37f48a;
mem[567] = 144'hfbc20bc700350a030d6cf52b008d04740e98;
mem[568] = 144'h0ccef026ff7b0dccfdf3f417f579039f05e3;
mem[569] = 144'h07a2fd25f31dffcb03aff561f551f2a10b3b;
mem[570] = 144'h01b1055ef9edf5d902b5fb85f8c106f4f713;
mem[571] = 144'hf8a4f96bfc980eb8f660ffc80361f7ad0350;
mem[572] = 144'h0924056104caf5ef048dfdcdfd22fb54fe1f;
mem[573] = 144'hf4d7f7e30ef005d40fd9f9adffbbf45b0f48;
mem[574] = 144'hfe2cf2650c700a26016bf17f08fb06a8f66c;
mem[575] = 144'hf2840892018e0466fa75f8c5ff4b0edef8a9;
mem[576] = 144'hf7950b21f26ff95000c6053a0ea4f69400eb;
mem[577] = 144'hf11f0b4002a9f6190c62f459f0e807fdf640;
mem[578] = 144'h02b9f94707b40040ef5c0976efc9094a0692;
mem[579] = 144'h03670b04f1a1056204ec059a0c7ef5b9fc99;
mem[580] = 144'hfd07f661f91eefc502290c5e0c9df8bdfdd2;
mem[581] = 144'hfe87058d0176efdff3fbf93309fb02460424;
mem[582] = 144'h07aff64bfcac07bdff8ff7faff9607870f25;
mem[583] = 144'hfec006970a7a0c3df925f5e3f30ef1acf5d2;
mem[584] = 144'h04fa05f2f3edfaecf4070a61f4aaf92706a7;
mem[585] = 144'hfd2d0c21f9640cb206a806860a37fa45f721;
mem[586] = 144'hfef2f5c80c4107be0025f62bfcc7f46805bf;
mem[587] = 144'hfeab02bc0f5c05590929f7a700940ec907c3;
mem[588] = 144'hf036efa902d60088072efefa038c0578ee8b;
mem[589] = 144'hffba0780f593fed2f6930b4506c0fbbf02e8;
mem[590] = 144'hfa33f7850ad10373ff21fc8e02f7f502f5b2;
mem[591] = 144'h03fc066ef25eff7707dff22f0caa0ea60e35;
mem[592] = 144'hfaff0abf0c8bfd71f113f2abffd7f15eff07;
mem[593] = 144'h06e5f38b0d0bfffc0a8ff5ee060706a40149;
mem[594] = 144'heb0cfaa70cbee895f48de7c0f1eb03860f2b;
mem[595] = 144'h05dd0a60f85ef35bfc4e09480654f09f0864;
mem[596] = 144'h0a52f864f516f9700335ef01f1690620f6f8;
mem[597] = 144'he97afcd3f6580b78e5f4f8120582e684093d;
mem[598] = 144'hf5950d8e00b5f91af2ce0b2df4fc0062075f;
mem[599] = 144'hfc750bc0f8a400800c4b0490f168fee6f793;
mem[600] = 144'h097cf8a1f83afd65f804ff90f83bf09b0637;
mem[601] = 144'hff7bf74608a8f343f2a1f5d2f66ff6b6f6be;
mem[602] = 144'h03fff7bcf2d7f1d504c7f0dafb7504810569;
mem[603] = 144'h0f39088d044e0ac1015d0de40c4e0babfe3a;
mem[604] = 144'h1923fe50ea40fc2ef692f9c409da0ffaec0d;
mem[605] = 144'h028bf432f22eefc1f706f0d2f7adeec304ce;
mem[606] = 144'he5aee3eff5b60cb6eeb3026be82401c70915;
mem[607] = 144'hf85dfcf7f9a9fe26f165f25105dcf597f104;
mem[608] = 144'h04d90238f092068ae38ce0b0ffdff54cfd47;
mem[609] = 144'hfc640161f7b106befd81fb70efd7f7c8f8fa;
mem[610] = 144'hef3dfa610246fe420725007d01a8f1fdfa61;
mem[611] = 144'hf4810819fae1f0f2f3edf059fa94f2d401a3;
mem[612] = 144'hfc01f656fceefc6df9500d2b09a80b9effc6;
mem[613] = 144'h076bfc70efdbfaeaf208f9f40788f122feca;
mem[614] = 144'h0a03f5410d750b1f0a230d38f527fb56ff33;
mem[615] = 144'h0bc6087d0acff7e5060f035ef541f2cff3df;
mem[616] = 144'h0a8dfe5bf305ff69048808dc062c083d0928;
mem[617] = 144'hfb15059306460a44f502f63bf449f417f28c;
mem[618] = 144'h0c21096df48bfb4a01fffd8a08a8f676fea1;
mem[619] = 144'h0e670cccf72b0a05efd2fd0ef32f066cf045;
mem[620] = 144'hf8c3030df1060a1205ee0574f44fff6102f6;
mem[621] = 144'hec4e02f4fdf30b52f78c09210860f93f0993;
mem[622] = 144'hfdb90b21f6d60504f12efc3c0ee207d7f378;
mem[623] = 144'hf692f25df464f7a3007e0b4cf2baefc3f5a9;
mem[624] = 144'hf00ef33cf5f60a05f93cf37407eced730d9a;
mem[625] = 144'h0cd30cc1014f0b4202fb0ba30a2a0caaf944;
mem[626] = 144'hf836fa910c8df955dd2bf1e8e49df650f6b0;
mem[627] = 144'hfc3ffe780882f2890623faa6fd66f8f8fc49;
mem[628] = 144'h04aaeecdff6efcd9f1100cbd0908ee65f78e;
mem[629] = 144'h0660f59105acf366eaa2e561f557e3d5effe;
mem[630] = 144'h041af5b50c73096a05b709a4f29a064dfac8;
mem[631] = 144'h05c3fab6f828fbbeef4efe5df973effc0c31;
mem[632] = 144'h0c8cfbbbf0ae0b84ff2df18f0495f52201c0;
mem[633] = 144'hf44a07b0f248081b0cb7f760fcb2f9740c86;
mem[634] = 144'hf0eaeadd047e0b6fff2f026f05c9fff3ef73;
mem[635] = 144'h04fd019cee6107d70656fb1c0040f4d0f0c6;
mem[636] = 144'h090bf61de293fec3f53dee1911b90962f40f;
mem[637] = 144'h030a0a11fc12ffacee65f684fe7ef8fef11e;
mem[638] = 144'hef4cf2cbebf7efeb078bf242ed1cfa93ed9d;
mem[639] = 144'hfe5bf5e9f4bcfb8bf29c091d0306f9bdf975;
mem[640] = 144'hfc01f9c4f939fcccea99e05df64a01fdf47d;
mem[641] = 144'h05f3efb4ff32fca90351eb2ff63df97afd87;
mem[642] = 144'hf9b90c28f18cefe8f85efe52ffa9f061fae8;
mem[643] = 144'h08460ad7f5ecf0540095093e04c50721007d;
mem[644] = 144'hf0faf61b0ad8fea20c200d4cfe7ff204f01f;
mem[645] = 144'hf79800edf387f994f6970281f4c6f783eea3;
mem[646] = 144'hf0fbfa880f79fa5e0194f643f4ee0302f81a;
mem[647] = 144'h04d9ffb105a8f827faaffeb30129f6af058f;
mem[648] = 144'h0dbd03d3fc270593fbe1f697f497fd8f0f1e;
mem[649] = 144'h00afff850d450110f839fb35f2c5f8b30a49;
mem[650] = 144'h08880271f4ca0c62f9d0f68df3650fa80677;
mem[651] = 144'h0cc70baa04db0a2ef676f99e00f1f78f0c0d;
mem[652] = 144'hf7d1f7ce0657fb170637ff6efd3600ef0352;
mem[653] = 144'h0b7407a0f12ef77108ae033b0a350c51f783;
mem[654] = 144'h05150b91009b0219070c03e406000b65f223;
mem[655] = 144'hfa5d03200ff4f538f573fb46fa60f53af73a;
mem[656] = 144'hff4d0530f1550e7df40e0482f832f94ef909;
mem[657] = 144'h098ffe3c0da504000285fe9005a8f2e6f0d7;
mem[658] = 144'hf8fbf86c0183f9e5f92afab6004aedc1f285;
mem[659] = 144'hf9250d74fc8df59ef29e0e31f86c0867fc25;
mem[660] = 144'hf515fe5708e9fe860a18052df36305160d87;
mem[661] = 144'hefe6f4a8f0c90d40029ffb2c01d20c3405dd;
mem[662] = 144'h047ffb130022f751f983f1a3f845fa7e027a;
mem[663] = 144'hf45403c9f003f3dcfcd0f01b09d6f5ecfa9a;
mem[664] = 144'h04510428075aff8efb7b0b13f08cfba70c95;
mem[665] = 144'hf885f9480a6ff43d0b4f0c0eef8ef20702b0;
mem[666] = 144'hf0840d3f087cff4601abf5a10814f804f291;
mem[667] = 144'h0eb1f8b9febe05d0f367fb12f9daffcefb15;
mem[668] = 144'hfc42f41af7a7ee350514008af8f0029a0874;
mem[669] = 144'h01540b07fc94f0aff2affe5defa8f7cc0aa2;
mem[670] = 144'hf7f00bf6f4070a64ff18f1b5fa3d0b8ffcf9;
mem[671] = 144'h0f0801eb03680e6f0586f18106a6fdf4f5c0;
mem[672] = 144'hf33ffac601720c84fd56f422f6a3f031f6db;
mem[673] = 144'h045ffbb30cf3f8a3fecef62d0d9dfb40fd75;
mem[674] = 144'hf54df7cef0180601085df0a30b0df0250435;
mem[675] = 144'h0ad7f0c60634f2400cd00fc8f48ef4bff225;
mem[676] = 144'hf2fb05cf02ac018afbee073cf29d01fbffcd;
mem[677] = 144'h0384f17d01220ef007de0ca005c5faa3ef97;
mem[678] = 144'hf236012b070dfe48fc47fa9efbfcf1a7f36a;
mem[679] = 144'hf46308affac5087a0f6a0c190e380236ff5f;
mem[680] = 144'hfc45f20e04fc0b9e0bd704020dad0147f1f0;
mem[681] = 144'hf83209f5f62a033c03d50b21f150f3f0fd20;
mem[682] = 144'h0f39f91bf101fb2af178f19900c00f33f715;
mem[683] = 144'h0bcffde10c75f27dffba00a5fa15053ffbe6;
mem[684] = 144'h0c5ffb540cdcf272075ff2760b81fae8006c;
mem[685] = 144'h013ffd550e350e6b0ab10cb2f3c6fa45fa95;
mem[686] = 144'h03be0fb60d9df63bf21cf486f1ca0b86f68c;
mem[687] = 144'h04f8f898f1e409cb0b52fb0100c4f18efd48;
mem[688] = 144'h03fd022efc70fbd2f89df0240b9af0fc0dbc;
mem[689] = 144'hf5850d5b04aff0ebf51e0e2300f4fd9ef062;
mem[690] = 144'hf65a0cdaf4710b2df83cf16302b3f4c5fbc8;
mem[691] = 144'h04b706cd0a4cf0cf0b41fc90f8ef091308a4;
mem[692] = 144'hf317fee2007800d2083af202f553f786f6e6;
mem[693] = 144'h08fffc25f495f242ff220317ee870c92f7e2;
mem[694] = 144'hf1d100f9f45906ec07500ae00370077a057f;
mem[695] = 144'hf9e20c8efe6102df083cf98e00aefd2dff9a;
mem[696] = 144'h0d7703980e8eff2d041d064e0776fc410809;
mem[697] = 144'h02620ae2fe770caff206000d01befe63f54c;
mem[698] = 144'hff1709e2fd27fa97f41efd2b0652061a0091;
mem[699] = 144'hf0cffea5f27ff689fc02f32307c404b0f3c7;
mem[700] = 144'h004decbc00b1f096fb49ef9200d9f1a40d66;
mem[701] = 144'h0b15f754fa1af31e08330abefdd201d1071a;
mem[702] = 144'hff050ae3fa49f720015eeffcf743f1680159;
mem[703] = 144'h000cf76c0e70fe87070ef5e402430f4bf392;
mem[704] = 144'h086bfda5fa29f4b4058cf2e6f41e07ecf0ce;
mem[705] = 144'hfd4ef0d9f8f60ccc014ff585fa91f5e6f98d;
mem[706] = 144'hf1f10d62fcf8ff7408240687f854f43c0c5c;
mem[707] = 144'hfa6dfec8016ff992f186fdc5fb12f5240857;
mem[708] = 144'hf5eaf418f98b0021fdd8f442072e0c800c4f;
mem[709] = 144'h0c37fb7aef590e7904befadc00d7f173005d;
mem[710] = 144'h002ff300f5b0f2a40555efb0fbb30f96f62b;
mem[711] = 144'hf010062df92cf69b012004560c0cf68cfbe1;
mem[712] = 144'hf6dfff8f0027f189fe53f3630306fda9001e;
mem[713] = 144'h059df8ddf950f7500a99f2f1f802007df226;
mem[714] = 144'hf510f430f4c308cb010ff713fad308150379;
mem[715] = 144'h08ed000f0e590903fae9f608f70d0d89081c;
mem[716] = 144'hf130f9d706a4f0400481f1a7fd85ff23fcc1;
mem[717] = 144'h0721f07e01a6f73a0427f0a0f170fe2d0a81;
mem[718] = 144'hfb250683f1d0014dffa6fda702450de4fea1;
mem[719] = 144'h092e064000f3f4bdf2ed05c0014900a707ed;
mem[720] = 144'h0210058cf9820e7d0d59f5f5f886f90e02d6;
mem[721] = 144'hfd7df4f90297fa64045f04c209960a460215;
mem[722] = 144'hf638f472f7160d14ea1ff22fe5e1ff47fd24;
mem[723] = 144'hfe7c02560cc6ff6f0282fa1cf2820671021e;
mem[724] = 144'hfdb808050535075afe0407a7fc88fc77f1f4;
mem[725] = 144'hfa00ece3f7eb024cf322ed77fa8bed64f03c;
mem[726] = 144'h0272fc4bf597074fef34f298fc1200a70b58;
mem[727] = 144'hffe800a605e7fdfd02640863096cfdd2fc2d;
mem[728] = 144'h07f9ef6b031f02b6efe10c32fb08f48af485;
mem[729] = 144'hfe9cf0df0241019b04fc00c2feb7f8d20b7a;
mem[730] = 144'heeb002c7fc420bdf08f4fbe00ea8f901fd59;
mem[731] = 144'h0ee6fffcf0e3fb2e01c0fd36fc900803f378;
mem[732] = 144'h0b98fdf6f257eb1efb9408bdfba90ab600f3;
mem[733] = 144'hf2d209af09e0fb22071e073d0105feeef784;
mem[734] = 144'hf562f4290866f3820d1a0783f2a6fbf8f08d;
mem[735] = 144'hf3ba03ed0d72fa390da10708fa03ffd3faa9;
mem[736] = 144'h00410155f34e01f0ff1d02e3f9b0f9b70836;
mem[737] = 144'h0197f3bff5480061f08deec9f8a400a4fe2c;
mem[738] = 144'hf59df23a010efd720ae20739f04efd250c56;
mem[739] = 144'h0a990f4e0d4cfc710c2bfde7f6c9f2580395;
mem[740] = 144'hf568f26c040ff92901c20ae20025035000fd;
mem[741] = 144'hfabc066b0385094ff888f31b0bcafdb8fdad;
mem[742] = 144'hf7f9fb380d27f85e02eef7c20715f56d0384;
mem[743] = 144'hfada0e83f448091bf2210bd3f31ef88f0caa;
mem[744] = 144'h0c6deffdfb12ffd7f7bd08e203a5f6dcf0ad;
mem[745] = 144'hf2a8fd92f74a0603021c017c02d80202f8fb;
mem[746] = 144'hf7bbf496f5700cc4f4fb070fffd7fc64013a;
mem[747] = 144'hf6b20f8201e306b6f6e0f9630d82f87ffaed;
mem[748] = 144'h089ef20bf3a903f005a9ee81f95eff27fa2b;
mem[749] = 144'h0c280bcbffd20b33f313fe54f7a6faabf802;
mem[750] = 144'h0951f02f03bb05b1fc69025d08e5f8c40fa9;
mem[751] = 144'h09aaf2a60c1cf5dfff350d740fd40c5e090d;
mem[752] = 144'h07d60763fa2afb31f37cf9f90c35f8020cfd;
mem[753] = 144'h0533090d090201ed099001090b3ef402f057;
mem[754] = 144'h081e08fcf9f8f8620d890733038602fef72c;
mem[755] = 144'hf7c60b1a03cb0fd8fb2008a301c9fc9a02d8;
mem[756] = 144'h00acf3f008d8019df7dbf34b0d70fa10f573;
mem[757] = 144'hf0010e89fc7a0dfffc1b0222f3140cfff44a;
mem[758] = 144'h0f790112f29cf41c05f6f422f829087df11c;
mem[759] = 144'h0e48f2830b4302c0057509a0fd0fff50fa20;
mem[760] = 144'hffa4ff95f7e00e0604f40532fcebf0de0f1e;
mem[761] = 144'h0473071f05d7f108f064f045f5acfaea0a60;
mem[762] = 144'hf1b0f116fcd9fc16fdf6f6d708ec0b770d1e;
mem[763] = 144'hf3dc0bd4f9d30957068e01dd0141f155f83c;
mem[764] = 144'hfedff37ef3570a61f522f00b0b130db1f729;
mem[765] = 144'hf31e0abefc90f524f81bf51e0159f0ccfbfa;
mem[766] = 144'h06f001c4f3f8f3f5066802fd0afefde00d18;
mem[767] = 144'hf5660724febafe2e0d000763f3d0097bf43a;
mem[768] = 144'hf822f2f60e65f3a9fef20b41f01ffeb60da7;
mem[769] = 144'h0025f87bf2500043ff2709ef08fbfe7a0ef1;
mem[770] = 144'hf91bf42306adff1df5c7f2050645f8d6097b;
mem[771] = 144'hf0950f400d22fe1105340816f19b0a1b03bb;
mem[772] = 144'h059a0bdc0bc50263f409081cf6dff4360ee0;
mem[773] = 144'h0cc8f142017ff261f98704bc02cdf36f0be6;
mem[774] = 144'h024d0826061e0e5e07fbf0fd05b30fa90b1e;
mem[775] = 144'h072af5f409320d35f0b9fb7af53705b806a5;
mem[776] = 144'hfb78098a0e6df02b000ff2b904ba0103f213;
mem[777] = 144'hfeb9fc1b072ffa5709980049f1c50a430b59;
mem[778] = 144'h0906f7e40dd90816f6880350f0baf32cf258;
mem[779] = 144'hf50cf414f377fd4df8a0f2ddf3e00b77ff56;
mem[780] = 144'h07fa06300abe0661f5fe06c8091ef4b3f1e4;
mem[781] = 144'h0d25fe1c023900c0f86806f808f70ca20ab3;
mem[782] = 144'hfd460acaf841f61afb6b0584f8e00834f129;
mem[783] = 144'hf6bd0379fcdd003dfa120021f36cf89f002b;
mem[784] = 144'h025904a4f17e0e9e0275efbdef23fde2f933;
mem[785] = 144'h09cff052f467f923f16a02e0f67c098dfd99;
mem[786] = 144'hfd4afea402bbf50cf1380efcf87d02490b6e;
mem[787] = 144'h036cfb090c99f4cdfe620fbdfd4e00f4f7ab;
mem[788] = 144'h0baa05e4f0d4f6800364fa42f4500db10e3e;
mem[789] = 144'h004807ecf1b50e52fc6f0271f3eaf36900ef;
mem[790] = 144'h0df0022ff5f10a0cf6f30c9ef10dfa58f45a;
mem[791] = 144'hf38207d905bc07f7017309760059f61d096c;
mem[792] = 144'hf7000672f5350ecffd200a0501da06e305ed;
mem[793] = 144'h0f9e08cbf286030c0e6cf8150e400b7100f7;
mem[794] = 144'hf5d6080cf930fe33061cfa76f7acfd38f5b2;
mem[795] = 144'hfba6f70deff4f0210e95ff0501300e190494;
mem[796] = 144'hf394072805e902a6f24cee9cf0f5f7710667;
mem[797] = 144'hfed80da7f382078400f0f129ff5af342f017;
mem[798] = 144'h05f7f3070276fd470fce0bd7ffdbf394f590;
mem[799] = 144'h04ce025effa6f7ad08bef47f08e10e53fb84;
mem[800] = 144'hff6806c1fd88f03300fcf875f4a4f971ff53;
mem[801] = 144'hf54bf4ee03bcf817f2b30b23f267fe27f456;
mem[802] = 144'hf186fdeaf79ef49401280750fd000282fd9c;
mem[803] = 144'h0128f8c8fb0208a9fe0cf64a06b00e360932;
mem[804] = 144'h082d005d03ad01930354f76cfe180ea5ffb6;
mem[805] = 144'hfa07f525ff86f752fdb20da5f613f9be020a;
mem[806] = 144'hf727f4de09ecf3bbf6c20e78fe170757f723;
mem[807] = 144'hf9e100cafc6a098f0f34f0d8f050f4b20ef7;
mem[808] = 144'hf70cf76400dd0a6808370f8df5fcefe50d3d;
mem[809] = 144'hfa9f04520259019b0871fe810556f82104d2;
mem[810] = 144'hfca40d17f46a05e1f7aff31b066f08ea0891;
mem[811] = 144'h0620fee7f2a80b7a068ff2740c40f22200a5;
mem[812] = 144'hfba40a20f78b0d22fbb5f096f5b3efd4fa63;
mem[813] = 144'hf6bdf025f1480af0fb980e5df9ccf6310001;
mem[814] = 144'hfe58f2690f770963f76af1e1f21f013e049e;
mem[815] = 144'hf5ef08c3f0c008620ae807d7f9fb056d0938;
mem[816] = 144'h0c3f026cf3290479f1a4fb7dfc7f062eff72;
mem[817] = 144'hf847f1cc0071fdd7f78ef4bcfd62fad9f28c;
mem[818] = 144'hf0ba0359f20cf83ff02bf044fba6f3e402d7;
mem[819] = 144'hf73efa200fe207b7f08bfc030c23fa220694;
mem[820] = 144'h0f7e03baf658f6daf7840adef71b0fa8f55a;
mem[821] = 144'h02acf019f2bcf6f2f7560806f0effe8000fb;
mem[822] = 144'h0b08f649fa610765f07afd9209800809fc04;
mem[823] = 144'h03990cde0bc00742f87cf68c090a0bff0105;
mem[824] = 144'hf803fcf70fe70828f808f536f2a3fc0a0773;
mem[825] = 144'hf75cf0dcf71af84efab9f703075af1270ec8;
mem[826] = 144'hf322f9970d3907e2f2b10a25fdf400aa0458;
mem[827] = 144'h0c82f3eb07e70f6ff01afed2fd1ef9100dcc;
mem[828] = 144'h008d0482f7a2078e02a205c406e3f170f7f6;
mem[829] = 144'h0f9af1ebff88fa25f2d702fdfbbbfbe3084f;
mem[830] = 144'h02f208690c700d12f302f6a501a60e14f1c6;
mem[831] = 144'h099ffad5f0100e2d0cb2f2c30eae09cb059a;
mem[832] = 144'hf156fd75040af61502c9fb25f03a0464fa3d;
mem[833] = 144'h043108a7fa1c0c1af539079607cc0a5605af;
mem[834] = 144'hf56cf3e1f00b07c60a2304f5f15cf233f2d0;
mem[835] = 144'h0d54fab70c71f2cb0b7e069902fa02750796;
mem[836] = 144'hf6880a870baa01780b1dfd5af766f71406b6;
mem[837] = 144'h0a64fafdf696f3380c9bf5490721ee760ab2;
mem[838] = 144'hfdf4f090093cf793022cf3f1012d072ff61c;
mem[839] = 144'hfe90ff0ef5b60ad8f9c904dc036f03ebfcb4;
mem[840] = 144'h004506530d0a080ef7e20cd40709f7160ad8;
mem[841] = 144'hf12cf1c9f29cf7b807360c1b015cfb1cfb3b;
mem[842] = 144'h08f4f0290d66f4bcf2a3f201ff05f485f47c;
mem[843] = 144'h0b3bf648f16afe7afb8701eefb6cf172f857;
mem[844] = 144'hfc1d088b0801f7f208c5fb4afdf0f14d0831;
mem[845] = 144'hf59bff15038901840609024700210528fbe3;
mem[846] = 144'hf8bd03540839fc7b0871fe3d0b2f021f046d;
mem[847] = 144'hfffcf024fdaffcb5f676f066f7ab0bdc07b8;
mem[848] = 144'h0b790d09f3c2075d01dcf2d3ef31072c05ef;
mem[849] = 144'hfb880e2307c40eaefd5e0674f51c08fa0543;
mem[850] = 144'hf69802fef5f903490c79fd2af1a3f0e8f7d9;
mem[851] = 144'h0dae017dfb84feda0df8f51bfe9af611f458;
mem[852] = 144'hf55af0480daaf21af3ab0518f8bdfbb1082f;
mem[853] = 144'hfbcbf1ebf48b00dd095b01f1f5f2fbb1ffcd;
mem[854] = 144'hf125ff2609e7f31606a00ec502ce0534053a;
mem[855] = 144'hf4f40ea4f6bb03470f2b02f6001b01da0acb;
mem[856] = 144'hf582f93904d5f5a2ff940343007f0d7a0998;
mem[857] = 144'hf08201b7f5e6fa710f74f61fff54fe5709c9;
mem[858] = 144'hfac70545f56b051d0f370391f55ff4ba03e6;
mem[859] = 144'hf9c9feddf5b30a5df25bfb4bf415f643036c;
mem[860] = 144'h06fd04e1eeb1ff2bf03d01f407ca0144f88e;
mem[861] = 144'hf6be0bad0b2cf4e1fb59f15cfc8ffe08f83b;
mem[862] = 144'h0b94f064f26df10c0b2bf5dff232feedfb76;
mem[863] = 144'h0d6e0ca104d904fa039af49e022cf39909d8;
mem[864] = 144'hf7e005f1f68dfcfa079d03fbf8210ad7f216;
mem[865] = 144'h04cdfbe1036df11eefeb00a607ccf57cf610;
mem[866] = 144'heee8f024ff7b06cbf8e6e9e5e646ec5f029d;
mem[867] = 144'hfed5f89208c5f8edfe1bf9a407e3fc09f007;
mem[868] = 144'h0c1b002d0af40aae0a1df006f431066ffe45;
mem[869] = 144'hf88ff377e77cf755078afb01f521e46800b4;
mem[870] = 144'hefb9f169f934f6770a10013b03ec0c8bf2f8;
mem[871] = 144'hf58ff6760dda033103d10948f1a90079f4a7;
mem[872] = 144'h03ff0beff41df9d40ea5f5700040fb7bf329;
mem[873] = 144'hf2dd0c720f4e0b7ef559033ffb6df9b704b7;
mem[874] = 144'h0c160dc9f07bf3ca0e8c0804f444f86af28c;
mem[875] = 144'h05be079bfa53fd7df83a03e90c79fcca05c7;
mem[876] = 144'h10b70226edccf0f009c7f665eb710a2df8b1;
mem[877] = 144'h0564f3020212fa1802f4fb98f057f5cb0c83;
mem[878] = 144'h0437f54af4210c52f99efd3ffd1ef142f695;
mem[879] = 144'hf4810d30f3eafa1c0777fb11f0000c480cb5;
mem[880] = 144'hf2b3e7a80432f826e932f461e90a00b6ebef;
mem[881] = 144'h08ba082103010169eeb5f5d7f765fb2b0405;
mem[882] = 144'hf9b3f32d03a1082ff5f0f1e204b0ffb2005d;
mem[883] = 144'h05f30d10fa51fca601e80982f9ae0fbd076b;
mem[884] = 144'h0c8ffc3cf139f661fc120776f53af0c60aba;
mem[885] = 144'h083bfe170a4f09f40887082afff808bc08dc;
mem[886] = 144'h07d7004cf60c08f7f0e5045c045dfc1f0a24;
mem[887] = 144'hf3f205dffdbaef4bf54cfca0f6e7fae2fed2;
mem[888] = 144'hf460f1a007170dcf06ca05bbf06a0bc506ae;
mem[889] = 144'hf566f3adefe1fe69f4f3f5bef10d050af713;
mem[890] = 144'hf55ef745fbdc05370b14ef0ff15bfa4a084b;
mem[891] = 144'h09d405c7f481ff0cf93cfcbff254003af62e;
mem[892] = 144'h0594fae000b5f1acfcd706c40390ece805a5;
mem[893] = 144'hff87f59700190344f9120763f93bf3ee0d42;
mem[894] = 144'h0279f0b7f9270a1ff5fcfbe50c4dfdd5feab;
mem[895] = 144'hf5b0fd510c98f21a080cf9b80a8a08e7fbf9;
mem[896] = 144'hef2ef5e10ab0f4a6f993fe70f726f92bfb18;
mem[897] = 144'hfc3d03bc0633f669090507c9efe60708fcbe;
mem[898] = 144'hf0aefd9af3cb014201c2f1e8f5770a8e0d06;
mem[899] = 144'h004a0560f4d2fdaf0fa9f6d3fbd6faf609e3;
mem[900] = 144'hfbe6f1d500ddf74bf8dc0f3bfb8402fc0aa8;
mem[901] = 144'hefdf0271efe2f269f5b3fd5eedeafe27f253;
mem[902] = 144'hf21dfb21f4a3f5f8fd3bfb9506b005f605c4;
mem[903] = 144'h0e6b02a202ee0196014f0bee0de207b4f545;
mem[904] = 144'hfd0803a9043df8caf42e061afe96f31f0f39;
mem[905] = 144'hfb290315f9f4f164fddf0464fad5f8c7eff0;
mem[906] = 144'h0133fb64081804ec07fdf7bb0ceffc9c0925;
mem[907] = 144'h035af2e1f106f63ef9a8049b08f2f657fc79;
mem[908] = 144'hf9cbfd0f0bdb0acbfa9505da0108091a0b17;
mem[909] = 144'hffba0d7506f10d7900ca0a96f21df93e09a2;
mem[910] = 144'hf800f41001b60683f77701430b7c08330074;
mem[911] = 144'h0dcb09d00519f078002e057bf60a04ea0a4b;
mem[912] = 144'hfd77fa07f4dcfadaefce024204690bbbfb36;
mem[913] = 144'h0594068a0b0bf5e7fb480127fcbdfa350da9;
mem[914] = 144'hf22ff808f3d4fe2a0dcc0263f6c4f93a04dd;
mem[915] = 144'hf8e508ec07710bb5fcaffa11f4210ce001e5;
mem[916] = 144'hf3f506d4fb88fbca0794fb680f43faff0223;
mem[917] = 144'hf52e0a40fdf1087502250a1a0b0c0a26fd1b;
mem[918] = 144'h0e1ffcc30ce30bca09150e59fae10b2bf91d;
mem[919] = 144'hfeceff4107cd0ad0fa81f2e0ff1ef0d1f679;
mem[920] = 144'h07e202a0093c0b4803880dc7ff9df053f2a5;
mem[921] = 144'h0b6bfaa305bb03cdf065f7c80725f6dbf346;
mem[922] = 144'hf3cf0731ffd5f025f3490e44f79cfbcdf863;
mem[923] = 144'hf929fb67f8fff8e4f37a037c0ad9f4ed09fb;
mem[924] = 144'hf87ff86e012006d4fda502c10338f7be05be;
mem[925] = 144'h03b3f747f18803aa0816fa18091df73cfcee;
mem[926] = 144'hf4cbefb10bd40f7fefee00d701580c750e7c;
mem[927] = 144'hfe2eff4ffe1909d409b70c00f609f4f108ab;
mem[928] = 144'h0e2c018f06cbf23b0b5af7e10b90f87df3a1;
mem[929] = 144'hf890fc83fa3201e3f270fefdef29f1d208fc;
mem[930] = 144'he73c03f0f9bcf55bffefe8ebdbdaeeabff68;
mem[931] = 144'hef8af4f9038805f4f626fd3c0399054ff138;
mem[932] = 144'hf3cd08c5f227f865f771ff4b0a4cfdd708ad;
mem[933] = 144'hede0e52dfaf80060f784f801f072e821f3ad;
mem[934] = 144'hfd68f6fd057005e9fdd90a5609f7eff306a7;
mem[935] = 144'h0daa04380571fd08efc2f461fe06fb09fd82;
mem[936] = 144'hf713084007c5ff700703f035f6bff04a0a38;
mem[937] = 144'hf2710889f7bf0d15f8f9fc25f37e0638ffd6;
mem[938] = 144'hf51cfb14ff2df8fe0b2803ee0e70fefa01ec;
mem[939] = 144'h058ffd43f31ef75b0dd60c430086069902e6;
mem[940] = 144'hed89e4b8ef55e776f98f0b4cec190300ec77;
mem[941] = 144'hf5600268efa00f20fbfd080e01bc00faffaa;
mem[942] = 144'h05ae089ef73708b3f943fbce0385fcadf147;
mem[943] = 144'hfaabf1e60202f75f0d1efeeef4b20de60297;
mem[944] = 144'hed54e9390b20f394ef0ee919eb9a0104fe8c;
mem[945] = 144'h019502920c2affdc0c32fd50f4a2fabc082a;
mem[946] = 144'h0bfdffc1f274068a0009f4230635efaa03ed;
mem[947] = 144'hf8a3f44b02f0eff90b51fb05f060f094fa1b;
mem[948] = 144'hefe206d7f7ed07ca007c090606eaf460ff34;
mem[949] = 144'h07130319f8f9eec2065ef108fba9fdf4097a;
mem[950] = 144'h06b3fabaf30a0a96fba2f41d0e35f51909cf;
mem[951] = 144'hf6150c1bfdf4f9830b4a0b33f82d0121ff1e;
mem[952] = 144'hf79e02bdf0d1f3e7fa8bf3530a65f4a9f8a1;
mem[953] = 144'h01a5010cf95903f9f9690e76ff8cfc5ffd6a;
mem[954] = 144'h042cfaa0049af39efcc8f8cb0c6b0d150d10;
mem[955] = 144'h0553f7590d19fca7088a0e5efc7d00cdffb5;
mem[956] = 144'hf578feb7faf3facbffff0af9f8b8f508009d;
mem[957] = 144'hfe910304f4a6f2baf74b0b50fee60af30b0c;
mem[958] = 144'hf04e0ea8f2cf0e2af235f535f223f94e08c4;
mem[959] = 144'hf6bdfb54003305f3f671f3f0f194f7baff3d;
mem[960] = 144'hef77093ff7c809750880f7c7ff0bfda6052b;
mem[961] = 144'hfbd1f8e203b204bbef71ff16fd21ffa203e3;
mem[962] = 144'hf95bfd00fd0df20e084b009c007a0d4bf2bb;
mem[963] = 144'h0517f1bef7a1f09f05abf231f6fcff5a0dd6;
mem[964] = 144'h0967f3bbf1defa20f724f51d02cff59e08d7;
mem[965] = 144'hfc7d0d49fc68ffdf09bc0b8f0b12f1eef07b;
mem[966] = 144'hfa15f8970403f027fd1ffc1cee9fefb1f7fc;
mem[967] = 144'h0e96f42e0388f1f2f662f941f8ba04e40f07;
mem[968] = 144'h08850b0100100371f9c3045a0db60489f188;
mem[969] = 144'h02b20ea3f92e06c001d4f25a094e06c9f751;
mem[970] = 144'h0e2d0842f4e902ad09e201bb047cf03bfac9;
mem[971] = 144'hf7b50309090cf14905befda5ffb5f0de013d;
mem[972] = 144'hf3e90a5cf70b072500aaee19ed4e0631f873;
mem[973] = 144'hfdd6fdebfee2f120f5a10a530e82f2cef525;
mem[974] = 144'hf654fc20f862f05b0d07f95af7a50000fa9c;
mem[975] = 144'hfd95f75df170f48e0c6600e2f8c8044205ff;
mem[976] = 144'h0724039707a9fe60f876f1dffaeefeb7fbc8;
mem[977] = 144'hefa9ef8f046407c7fe80f68d090e075701cf;
mem[978] = 144'h0287f938f8eef26707540d120049f6d3f138;
mem[979] = 144'hf4cd03c0f901f77ff55700100eff05960b47;
mem[980] = 144'h0a3dfa51f764f365f1a90cc4f79302a10ca3;
mem[981] = 144'hf3410dc80823f5fff94ced1dfb55fa96015c;
mem[982] = 144'hf12e0b0bf476f6b9fae9fbbcffe40ae50032;
mem[983] = 144'h0955f6b7f50d0bf9eff7f55a0caa01350474;
mem[984] = 144'h0064f501fbfd0723f72a08b10f6e091b0161;
mem[985] = 144'hfc4204600228f10bfcad081efecefe5e08dd;
mem[986] = 144'h07b4079e06510382f284f7d4032e00f70226;
mem[987] = 144'hf8eb0cc1f2bdf5e700d60f0efbf8f40eff99;
mem[988] = 144'hf8e5f1bdffb60a2c09c20313ea78ed10f5b7;
mem[989] = 144'hf6a90280f2e4f09cfe4105430b7fffcc0658;
mem[990] = 144'hf7530526fc12f342fdcef04b06600c10fe3d;
mem[991] = 144'hf255f1d50f2409e50f14f53b0fd2f8640e72;
mem[992] = 144'h014f08d003ea0cdbfc4ef8200a48f4090ee2;
mem[993] = 144'hf6c3f2bc0b6e0699f4b8fbd607290061feed;
mem[994] = 144'hfb01fea90405075a016f01e20723038907c1;
mem[995] = 144'hf6fc02a5095b0304f00ff8240dfffcb805ed;
mem[996] = 144'h0d3b0bab0de409a00a46f969f7b0fd480e78;
mem[997] = 144'h09b6fc5208fb023e093df36a0c82fcf6fa8a;
mem[998] = 144'h092b03f4f222fcb2011f0c9c06130192efec;
mem[999] = 144'hf3f908320493fdd9f39ef70b08bcfc750e8f;
mem[1000] = 144'h0dcb0e360c83027af579f1020482fb45095f;
mem[1001] = 144'hf397f580fd2afe7305000e4afa1cf239013e;
mem[1002] = 144'h0e42f16601c10901f929f1100127ffa00793;
mem[1003] = 144'h09a100420b74f4ea08f900780e68f1c90a92;
mem[1004] = 144'h097e01ddf2c10a7cf0ea02c4002bfa52046e;
mem[1005] = 144'h03440cca0457f7150354fb47f3ea0df1fb36;
mem[1006] = 144'hfd7f0699f4eff704fbca0dcf031b08a000ae;
mem[1007] = 144'h08e005b306b4f92500430701f9d3fffb0d26;
mem[1008] = 144'h05edf9de0bf6f56a0577fe8309eb09470b38;
mem[1009] = 144'hf0f407870bce014d0c9df810f4b60d3a0d52;
mem[1010] = 144'h0e4b08c5f6f1fae8ee4405a50a2cf670fa38;
mem[1011] = 144'h0c05fbf902af0d88f565021a0f50f4cbf548;
mem[1012] = 144'hfb1a059709d0f803f3a305b6f096f9a4f431;
mem[1013] = 144'heebdf989f8e3fe8b061302e0f52af96bf83a;
mem[1014] = 144'hf79607e407d0fcf4016cfc570d5cf28607b1;
mem[1015] = 144'h0921f86ff7de0c5df79a00f40a3df8fa088b;
mem[1016] = 144'hff330511f5be0526f0e805c7f7b5fe500125;
mem[1017] = 144'h0b4bf27700c6f936fd86f37e091d023f0f84;
mem[1018] = 144'h033ef9170a8606a4faa6f5cef785fc5e09dd;
mem[1019] = 144'hfc090cec00a9f28b0048022ff8490be4fd83;
mem[1020] = 144'hff3e09640d3cf38a012408fcedc306bffbe5;
mem[1021] = 144'hfa1f04cc0c3cf6cc0006f717f232f0640867;
mem[1022] = 144'hf3f00c33f632f67605ef056ff6ce08020b8f;
mem[1023] = 144'h043f054ffbdbf1ae08160b17ff9809ff09d5;
mem[1024] = 144'hf426f55d0aac08db0af1f90afc32efac0774;
mem[1025] = 144'hfc0e0063fb82054af0fa090e056f0d3208b7;
mem[1026] = 144'h075af53304b10199f695f74afc16f78af1de;
mem[1027] = 144'h02eef09df989fa39f5f6f0c7f1e401be05b3;
mem[1028] = 144'hfe7df7a2f136ffc300b4fea409f3fe7c0407;
mem[1029] = 144'hfa2a0e06f6a4056704caf4e108270c84017a;
mem[1030] = 144'hf129094ff5fdf6c7f4f80930f082fd1a0ec8;
mem[1031] = 144'hfb9b0650ffe20011fafbf1a30d2605f00be2;
mem[1032] = 144'hfa7c0b75f2f80b84f398fce0ff37fbdff612;
mem[1033] = 144'h06eaf34d0c540e5f0d440560f2cafd71fe7e;
mem[1034] = 144'h02410a00085a0dc9f754fbf7f9c1f0040cc0;
mem[1035] = 144'hfb4f0a6afb43f8b7f61a07d400380a6f0249;
mem[1036] = 144'h07bfff05f10905ab06670545f169fa3c0abf;
mem[1037] = 144'h0641f1d3f512faeff7c6078e03fa054e0323;
mem[1038] = 144'hfcbcf9bbf35606b80496f9070f7d091f0780;
mem[1039] = 144'hfef6f04bffae08830328013ff67c0d5606c8;
mem[1040] = 144'h0d15fbc908f0f110f7af0d080483043af777;
mem[1041] = 144'hfdba09a20ebafa4709a5fa80f57e03400729;
mem[1042] = 144'h0bb3f000f5e3f97dfda4f62cf3cb06fd0d30;
mem[1043] = 144'h0481f4f7f914fe230cba0361f5ca0e51f25b;
mem[1044] = 144'h0416f0b10ef5f13603e804d70699fcd907e8;
mem[1045] = 144'h0aa6fe7bfb5ef756f6b804ea09810600f34f;
mem[1046] = 144'hf1200956ef820b6904aaeeb80c3ef10d0ec6;
mem[1047] = 144'hfee501a901fffe180d86059107600850f0a7;
mem[1048] = 144'h0743f339fcd1ffd709b0085303f10c6ef992;
mem[1049] = 144'h05a30e43f0c1fd4dff7903d30a0e04cefc15;
mem[1050] = 144'h087ff020f0a4ff4008600d30fd790e920c1d;
mem[1051] = 144'hf691f7f4ff85f27cff5ff144fe15ff9d0dfc;
mem[1052] = 144'hefb306960c62f60af856f145f2f8fc5afd49;
mem[1053] = 144'hfc7bfdd3f225004bfb5af7a5f648016d09ec;
mem[1054] = 144'hf650072bf00b0899f7e3f8bf0e6f0958081e;
mem[1055] = 144'hf652fae10d6305fe07c2fe620260f52cf968;
mem[1056] = 144'hf23d0453fd09f819f71ff06b045c03fe0023;
mem[1057] = 144'hf589010af20a0eb50814f4ac0b20fab0f793;
mem[1058] = 144'hfcdd068bf2e806a2fa37ead6f2bcf4b6f183;
mem[1059] = 144'hf1f2ffc2f6fcf30505f3fd56fd320e6501da;
mem[1060] = 144'h04c2f8280da7034aee0a040606f30bf9f5e4;
mem[1061] = 144'hfdc1f483f2f20d56f221fd8b0579fe81f27d;
mem[1062] = 144'h0506faa0f001f25d0282ffdc0082f48b046a;
mem[1063] = 144'hf3c60b6006b6ef4cee8d02be05120abe0d5c;
mem[1064] = 144'h02ab07ed05bcf936f3fafa48f1060d7702f1;
mem[1065] = 144'hf5a00d8dfd21f0af05c8f86a01b9f75b088b;
mem[1066] = 144'hfade066ffdd500b7fe8bf3a2fde10bc1090a;
mem[1067] = 144'hf90c0d7bf76d06dbf2aff148f4830a5ef9d5;
mem[1068] = 144'h0801ef3a02b60c92e29afe3203d1e74e049e;
mem[1069] = 144'h0db0f6ebfd3c0d190897ee540d00f1ad0894;
mem[1070] = 144'h0480f446f177f3c7012ef0810696ff4e0a7d;
mem[1071] = 144'hf1660e3b00a0ff8bf1cd00830901ffbe094a;
mem[1072] = 144'heb3df141fd0f06baff7b006e021c05e2063f;
mem[1073] = 144'hfc32028cf92f0b09f729f5b7efa2fbf2f958;
mem[1074] = 144'h040c02950d5dfad7083d024a04c60a05f21e;
mem[1075] = 144'hf692091a0023067cf3f1046600820f9cfe99;
mem[1076] = 144'h0f1907cff172fc2df514f7b2f95ffd70fe2f;
mem[1077] = 144'h0148f91706940523f6ec03ebf72d09bf0c3b;
mem[1078] = 144'hfc0df04bfc99049107ec0503f271f368fd09;
mem[1079] = 144'h03ce02a6fa64f7ccfa300353eea8044df781;
mem[1080] = 144'h03c7ffb607fb0feb0eebf63cf2a5f6f1059f;
mem[1081] = 144'h0dbc0b20f3700394f48a0399fa3e067e0f18;
mem[1082] = 144'h082903d0f934fec5f87ff11700bc06a40ead;
mem[1083] = 144'h061cf7680253f555f45dfd41007effbef3c3;
mem[1084] = 144'hefdefc07f98f0a84ed6805fc014108b8ed91;
mem[1085] = 144'hfbc600ccf697f5750d82f85f00210c51fdda;
mem[1086] = 144'hfd75fb87f7f6012104e906faf6d3f9b909f3;
mem[1087] = 144'hfdd5f7ab04330cb30631f59d03e00fe9f75f;
mem[1088] = 144'h091303010adff8faf9f70b68f8d4fc4b098c;
mem[1089] = 144'hfa0f027e010309890985f2600d6afe35faaa;
mem[1090] = 144'hfc97ffb4fc14f11b0b9533f3020b0049f159;
mem[1091] = 144'hfc9ff78ff5c0045dffbffa180915f557f03a;
mem[1092] = 144'hfedffda50180eb61e910ec98f7cdf2400d63;
mem[1093] = 144'h00aeff520e03fd80f4a3f160ff5100f90588;
mem[1094] = 144'hfb4e0272f606f2ebf038f5c6ef2101de049e;
mem[1095] = 144'hf62ffa67f869f27df5d7e3460a83099b0732;
mem[1096] = 144'hfba4f247efcc007df072fa5f0b03efccf5af;
mem[1097] = 144'hefcffa430e2d04f0fbddf5f201b3f25a050e;
mem[1098] = 144'hfaa6f088f4efef84fda5f168fef90ce5efc4;
mem[1099] = 144'h028b07510210ffbdfea6f75e01cb06750d19;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule