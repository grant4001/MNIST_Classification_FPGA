`timescale 1ns/1ns

module wt_mem3 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'hfb180516efba03c9efccefb1f395f5bd0589;
mem[1] = 144'hf83ff87a00fff14dfe81f6140545f1290049;
mem[2] = 144'hf919ee7604f10754f2ab0291edda03a5fd7e;
mem[3] = 144'hef84fe18fb870b0c00160b760576f697ff76;
mem[4] = 144'hfbfbef9ff99dfadcf0cb08150756f27707e6;
mem[5] = 144'hf8670b8ff31bffbf0a7bfe01f01a086fee9d;
mem[6] = 144'hef23fdd9028ff42ef372f4d5051ff93806a4;
mem[7] = 144'hf23f09e6032b0012fe4e0546ff73fb77ff2e;
mem[8] = 144'h04500a2009c300860deb02000884ee710dce;
mem[9] = 144'h00d00b7ff098ff8704cd0a72ef8104e50c39;
mem[10] = 144'hf623fe29f84ef25ff17df7adf7ce0e0ef061;
mem[11] = 144'h00f8f5fef555070cf156facdf9620715fef6;
mem[12] = 144'hf46c0c44f8baf5f905a4f3b4f165005a01d7;
mem[13] = 144'hfe9efb8ff61ff8d9fadaee1afe58f2670a77;
mem[14] = 144'h089dffc0f4d9faa4fe7cfbb601b1f677f4e0;
mem[15] = 144'hf95cf531fe29034af5ce027004af0313f564;
mem[16] = 144'h00fc0327027cf5e1010fef39f4560009f8de;
mem[17] = 144'hfb6d03d4fa850a58f863f36b0187fa56044f;
mem[18] = 144'h04a30283f9a208e30219f614f687f18e0413;
mem[19] = 144'h09dd07d9fd8bf0e1fcff0377f2cffa99fb79;
mem[20] = 144'hfd77fea0f0bef5bc00060252f0ee05dafe51;
mem[21] = 144'h016ffd7bf497024df2b5f7920161057d08db;
mem[22] = 144'h03e0ef33024f085bfb6503c60c4fff79026c;
mem[23] = 144'h04f30485f72ff6c0efeefcf8fb85f0bd0bb1;
mem[24] = 144'hf2efeeb80016fa800b36f32c05ce0606fd0d;
mem[25] = 144'hf6f2ef6a0961ef73fb5d0089f369ee5aed08;
mem[26] = 144'h0b80f90408d2f4a2fbc102e50641f34805e0;
mem[27] = 144'h0c80ff7ef7d3fb96f580f1f6ededf53506a8;
mem[28] = 144'h026b093dfd360e120383fa6af47cf5c00186;
mem[29] = 144'hf27f00b003ceeffe0d44ff3b02640662f6c5;
mem[30] = 144'h028c097bf27c04b5ecc70976efaaf536eddc;
mem[31] = 144'hfd6cedcaf6eef1a3f4d9f36407d4085ced99;
mem[32] = 144'h0c71002c0686ef48f327fd77f6c6022c02ab;
mem[33] = 144'h07ed096100a40224fdc8053beecfff2d085e;
mem[34] = 144'hf35df1ef05e6ff8fec89fb5efe3305e7ef90;
mem[35] = 144'hf3d40893017dee13f1d504caed8b05d307ed;
mem[36] = 144'h080eef05ff24f1600b4ff33009e30ba7f411;
mem[37] = 144'h0bb8013b08cc07fcfa0becce0d0afdfcf2f2;
mem[38] = 144'hf5d6efd2f99e000cf108f0b5f6c2ef62fb81;
mem[39] = 144'h09b4f828f9d1fec604b00ba1f9eaece4fe2d;
mem[40] = 144'hffe9f33ffdc4086afcbf014a0683fa20f2f4;
mem[41] = 144'h0cccfe3cf102f19002430a1c0ae9f824f2cf;
mem[42] = 144'h0c13f669f908fdc1050b054df5c10cedf1ac;
mem[43] = 144'h0df50c8cec3d00b5099b00dff737f45607e6;
mem[44] = 144'hee07fc45f998fb7a0b32fa87ed7ff4f1080f;
mem[45] = 144'hee32f41ff9c008ceffb3ffcbeecfedfa06c7;
mem[46] = 144'h0134fa62fdcdfb48fbf9fec70358fa760bcf;
mem[47] = 144'hfff10490f99af819f52c0a28fe7f0266f2a2;
mem[48] = 144'hef3cf431fa96f8290111f53cf59fff980a74;
mem[49] = 144'hedd1f8790397f121f8d30b8109a40c15f456;
mem[50] = 144'heff00296055ff48a0bdb092af8a5f39afc79;
mem[51] = 144'hf60d093a09a109a4f9a8fbbd0883fa7b0044;
mem[52] = 144'hf43df52109b1ed6c08880ce0fa5efe540147;
mem[53] = 144'heff1f285fb25eecef40907aa01d00452eed7;
mem[54] = 144'hff710969f206097a0aaefe9f0b5505bef37a;
mem[55] = 144'hffe10bfd025ef16d0d0bf097eec3f871f418;
mem[56] = 144'h0d360444fae20ef902b2feaff292fe5e04c5;
mem[57] = 144'h044af27bf4e70004fe1e0330097501d0f119;
mem[58] = 144'hfb31f3970b390abf04c1075df89bf5e1fcdb;
mem[59] = 144'hf6fffe3207bb095b0d9e01b4fc4b0e510c93;
mem[60] = 144'h019107b5f22c0cedfc5601af0042fee20ca3;
mem[61] = 144'hf4260784fa97ee40f8bdf9d90874f06c0211;
mem[62] = 144'h0287f98d044eede0eeca0b8f0515fb500de7;
mem[63] = 144'h0427fce5ee4800c8fb59fab90280fd8e0d12;
mem[64] = 144'h0560fdf700ad07ecfb600bbdf5e9f25af06c;
mem[65] = 144'h0883ff99f2de08b0fed8ed05f8ee090a0881;
mem[66] = 144'h08e3f4cc0d5cff3c09a0f148fd4e05ce0647;
mem[67] = 144'h0c63fc1e004b0929fb350eb6f7a0fe880e5f;
mem[68] = 144'hf97202d5f56a08c80079f933f7f4060903c6;
mem[69] = 144'h08bef9a70d6d04d7014c02b30814fc8f0fc0;
mem[70] = 144'hfb5509e10dfefb2b0be5f32bfe9cf8f801fc;
mem[71] = 144'hf21bfc24f27d0c45fba9f2a304ddf9d5f999;
mem[72] = 144'hf3ac08a5f6baf4eaf4170306f78a0a6af784;
mem[73] = 144'h0b2e0acef981f6510924f8cb0b63f5c4fb70;
mem[74] = 144'h02bd0bdbf776029902aa04bd0740fe2bf18c;
mem[75] = 144'hfdeafef40c5bf3a00f2cfd1ffddcf69df1ca;
mem[76] = 144'hf7f4f153000f0d08fb99f004f887f54e08a1;
mem[77] = 144'h0409f927f10c085c0beaf1260208f28efb13;
mem[78] = 144'hfeaff7b50ae70b840ec202f404dafa780f9a;
mem[79] = 144'hf8c503a603bbf11c03a2f286f41ef30af444;
mem[80] = 144'hf7cb065d0375010e0725f4f2fbc0f074f123;
mem[81] = 144'hf6380c01fa8d0e770690035df8560f8ef9c8;
mem[82] = 144'hfda7faadfdbf0fd6f996002607ac04d3f30c;
mem[83] = 144'h062e0879fa8a033e0c16f8a304ea0387f054;
mem[84] = 144'h0106f533f8c6004902790bc1f83af7dff24a;
mem[85] = 144'hfe8b0e46058201a6fa4efa220b200c97fa12;
mem[86] = 144'h0f9ef67205e6febef1bbfbcd0baa0a24fa2f;
mem[87] = 144'h004c0fa6f24cf0e4f128ff49f63ffda500bc;
mem[88] = 144'hf87d00080e3af9c7f3e70b5ef479fe070c44;
mem[89] = 144'hfc6efc79fc30044303860f06fc95f72cfeb5;
mem[90] = 144'h00c6087a00aefdee068b03b8f106fa9507f5;
mem[91] = 144'hf4ae0e6bf3970f270d6b0e69fa370289f25b;
mem[92] = 144'h07fa0f380409083ef95d007ef41b0ab504f6;
mem[93] = 144'h00f1ff98f061f76af65408c9f594fd09f5e3;
mem[94] = 144'hf195f3340ee6fabbf793f4820edf0614f679;
mem[95] = 144'h01950007f1d60b1aff0ff0aaf3960198f858;
mem[96] = 144'h05390eb2ff260948f516f53f0c14f85c0de6;
mem[97] = 144'hfeecfc9dfd480887f244fe77ff26fc8b03f3;
mem[98] = 144'hf8f501b7f28dffb208ca0c9e0c93f798f7de;
mem[99] = 144'h0e0b0d2df00a0e4df0320e60fb890151f55b;
mem[100] = 144'h003ef5a2f028f0d2f0260b7ef6b6f883f607;
mem[101] = 144'hf7330882fd880088f7d1068ef520fee5f121;
mem[102] = 144'hfee506dd0592fd1bf247001908bc02d00fab;
mem[103] = 144'h017903bff0b00400f95808ac08c6fc3103eb;
mem[104] = 144'h07e2fa7701190787faddf34609b4f1b7f103;
mem[105] = 144'h05be03d60329f370023bf87e06030e6cf812;
mem[106] = 144'h07d6ffcffc34068b0053f6fd013af4c700cd;
mem[107] = 144'h02a8001b0b6a0a0af0670d6d03b20a860b9f;
mem[108] = 144'hfad1fcacffc5f2680a87f78201f5013c07a3;
mem[109] = 144'hfd510c07f6450b3e02590d85fe69f7fe0cd3;
mem[110] = 144'hf275fd880df0f295fde50b730e3affe8ff4f;
mem[111] = 144'h048201a7015bff08046405590f26fb2f0d23;
mem[112] = 144'hf966064506460e640dd1f4edf2790eb00803;
mem[113] = 144'h06ddf870efef0ab500b9fa18f72d0bb8f74d;
mem[114] = 144'hfaa60180024f001c01b0fc56f0d3ff460de8;
mem[115] = 144'hfd1e061d0294043206490cd0ff570079080c;
mem[116] = 144'hfff807ecfcb80f37fb45019e0294f439fabc;
mem[117] = 144'h0dd90a42fa2dfcc3f08ef22bfd870384fae5;
mem[118] = 144'h0e1505fdfc060e19f60cfa45fadafc71f0ac;
mem[119] = 144'hf9effce9024ff74b0afff4abf1fe03ddefff;
mem[120] = 144'h03580a9a0adb0313fc5b01a609a4f6e40724;
mem[121] = 144'hfee10a07f7220ef3f016fccd0f45f40ffae9;
mem[122] = 144'hf4a2030bf8f704cb026d0f9401010bfaf747;
mem[123] = 144'h0fbc0634f64c035403fd0e97064af1250ba4;
mem[124] = 144'h070ffd0bfa970d5bf5c5efe10f320601fef3;
mem[125] = 144'h0561f779fb87ff0bfcb70496ffc707d6024a;
mem[126] = 144'h0825020a038008eaf97b061c080f0d35f171;
mem[127] = 144'hf16900710230f70bf5590f3ff314f9600285;
mem[128] = 144'hfbfdf4d005a7f64800a10c9d0a80f4f302b0;
mem[129] = 144'h00ef0616f4aa0ae6f221f283f4a9f4b7f251;
mem[130] = 144'hfbb5f5220a9d0899019cf92ff4660de3ff55;
mem[131] = 144'h0a1c0f0ef5480c1ffad1f63afcc8f9220aad;
mem[132] = 144'h0d2a0e3ff0d9f7c1016cfea10ab9fb03f9f4;
mem[133] = 144'h03ebf39d0f8a014cf576f2e3097ff4300a8f;
mem[134] = 144'hf37ef5430b9a0e5601660cae07dcf395f8b4;
mem[135] = 144'hfb9bf75ffa4206ceff29f9b5f0e5090b08c9;
mem[136] = 144'hfad307500ec302ecf894f9ab05670c2ef93b;
mem[137] = 144'hf4be0e8701aa0e2f034af88e0d52fb330cc8;
mem[138] = 144'h094ff1ff010ef3ff0ee605eaf26502570992;
mem[139] = 144'hf2b90938fdfbf9070e91fa01f458f68d0491;
mem[140] = 144'h08980771efdb06d009dbfc4ff1e7078a00bd;
mem[141] = 144'hf94006e9f4a404a8fd4a0419fd350f8bf74a;
mem[142] = 144'h04c9fe140d5501350eccfccaf1eef712fc7d;
mem[143] = 144'h0dbc0345f179f0dffe590b5b0346fbf9f15a;
mem[144] = 144'hf623fe38055cfc1ef9c9f46cfd1d0c090486;
mem[145] = 144'hfc86fb8efea40fc0026f0da5f73efdfa0dd8;
mem[146] = 144'h096ef3bffb1dfc6b0761f77dfd92f7b70c3d;
mem[147] = 144'h09c1f402f63cf3edf9c2077cfaae0c200363;
mem[148] = 144'h075e050e0b590cd5f2f20b330b480823fd72;
mem[149] = 144'h0767f66d0822f8c10e6ef5e7f69a0ab30a4b;
mem[150] = 144'hfa2b0b0701d3feba0170066c03f90fd5000d;
mem[151] = 144'h07ee0edb00c1f26d005a0f730fe30302f6c7;
mem[152] = 144'hfb21f1120f970d2cf1240df7fd5a020e0361;
mem[153] = 144'hf7a1ffd0fa57049af7ef08f7007e0d720b6f;
mem[154] = 144'hf53df6e70467fcfef4b704480f850fd5fa5e;
mem[155] = 144'h02e8f4620fab07670cba00530f74010004a7;
mem[156] = 144'h0fcef7e30ad705a309f8f2a50824017afb38;
mem[157] = 144'hf1adf9eaf536f7d8f60902540aa0f88ff04f;
mem[158] = 144'h02bbfd7a07cf023efab709fc0445f3c4fa63;
mem[159] = 144'hf54bf1c40396f348fbc0f7f40a7601fff7cd;
mem[160] = 144'h0f6802bf07980b1e0c71f6b20dc1fbddf5eb;
mem[161] = 144'h07ba086df2c108ca085afd9a0e22f98bf8c7;
mem[162] = 144'hf13afcc008f3fe8108c1f66b0877f6b008ec;
mem[163] = 144'hfb6104a8f4a70a0804bdf598f88c0de10083;
mem[164] = 144'h0cca0167f68efe59f8b6fb21049a0c74f2ce;
mem[165] = 144'h0aa402c1fa31f4ecfa9cf5ef04cbfe18fa50;
mem[166] = 144'hfc64ff04f978fbcaf827f3a00714eff3fba2;
mem[167] = 144'h098ef472fca70edbf6a0fc7205f8049ef64d;
mem[168] = 144'hff090952fb910017fbfefd32fb4bf5f10888;
mem[169] = 144'hf6c20ac806aefd82f9a20680040dfc720259;
mem[170] = 144'hf6cff551f673f05e08cdfd94f102f88609e8;
mem[171] = 144'h0efef9f20508f0e408bdf1aa0f9e0143fb2c;
mem[172] = 144'hfa0cf7c2fef1013906d10055f9ab02310da1;
mem[173] = 144'hf3f20676f1da0692061a039e0291fce60495;
mem[174] = 144'h0e6508c1fe200411ff2109bafdfb0058048e;
mem[175] = 144'hfb60f96902bdf28e0d29fa8bf1a307d70755;
mem[176] = 144'hf18bf8d6f5e8042708d30120f94df8bcf622;
mem[177] = 144'hfcb9fa96f1f0fc6d0c4e00fdf49e0c03f3b1;
mem[178] = 144'h073e0a6806a8f4400cd3fc2b00bef8b8f094;
mem[179] = 144'h0d38fc2600280f480d7af359088009b60e10;
mem[180] = 144'h09c1031f0b87f1fe02dff7980f8506bb01ea;
mem[181] = 144'h02e5f020fc080c28ffe1f4f6f9340d450d23;
mem[182] = 144'h0a66067f0af4faabf69a0fbf054ef7d6f6de;
mem[183] = 144'h02fcfc9e0409fcd10d76052e0e4402b7093e;
mem[184] = 144'hfb5e07fb00ad094201ddf0c2f388f2510e1f;
mem[185] = 144'h027d0147f5620aac0676082dfc0b0be1f0ec;
mem[186] = 144'hf09cf152febdf5e3060a0ae2055bf7560fec;
mem[187] = 144'h0cb60d9af5e807d8fda203d6083a0f7bf214;
mem[188] = 144'hff2703c60e660f940e1900c2f1bdfce5feaa;
mem[189] = 144'h04baf1b9fb3c03be0673f278fe46f6d606ef;
mem[190] = 144'hf5e50dbdf308f7a5fe9c011901600216fc08;
mem[191] = 144'hf8d20a35f3be05c1021b00ccf635043dfffa;
mem[192] = 144'hf901f450f972fa5f0387084bf9e805a70075;
mem[193] = 144'hf914fbd8f92bf49c0c64f7c10004fad1f914;
mem[194] = 144'h0bebf5ea02e80845f46b0308082408d308a7;
mem[195] = 144'hf92c01f7f082f7660c94fa0cf7b00efa07af;
mem[196] = 144'hfe55f781f1cbf32df025f1a10f53f7e3055d;
mem[197] = 144'hfc84f8890205f5fcfbc3f89605cd08860411;
mem[198] = 144'hf4f2f95208e8ff9907710e08ff580544fc36;
mem[199] = 144'hf95b00eb04170a79f52508860c3bf4e7f879;
mem[200] = 144'h072f060704b409b3f938f75ff2aef5e8f80b;
mem[201] = 144'hfa2d03160cb3f482ffabf75af2c00311f8a1;
mem[202] = 144'h0818014bf35d0887f3c40e9bfd10002a0be2;
mem[203] = 144'hf89507230f400e0d06bff834fb340fcffa4b;
mem[204] = 144'hf6960c4e02baf3fb08610c94ff88fb1d0189;
mem[205] = 144'hfafb0e800f6f0e0c0c69f5bdf7fb0923f9ee;
mem[206] = 144'hf031fb8bfc0c025506fef262f8eb016705d6;
mem[207] = 144'h0561fc6506e10175f323feab031809cb076b;
mem[208] = 144'h0e4c0673fa2607070886fc520f210ca40267;
mem[209] = 144'h0907f4e2f429f8c6054001b1009ffdfcf0a3;
mem[210] = 144'hf91f0001fc0a02150966f88ff569fa9405ed;
mem[211] = 144'hf522f643feef0d350fe7fb220eaf00b80668;
mem[212] = 144'hf7850a3bf727fbc6f0f6f44d05d8fe71f3b0;
mem[213] = 144'h039904f7074efde50503f5b1f9bff6cff243;
mem[214] = 144'hf726f7080ee40b35fcd408f6022203bf09b1;
mem[215] = 144'h0590f313fac9f902f8fe03740e98f1360a7d;
mem[216] = 144'hff85ffdcf4ba04c5f08b07ccf5d90ec3fd3a;
mem[217] = 144'hf0a4fe0ef1cef5300ed1fd85f74b00aa0807;
mem[218] = 144'hfd360e54fb4df47908440e8dfb59fe3efa7d;
mem[219] = 144'h04750bcc019200adf247f9e506cdf85f0ea2;
mem[220] = 144'h0905f786f8250c8004c1fdca0f50f5fbf025;
mem[221] = 144'h07e9ff1e076af55ff4fdfb22fd8b00f1028f;
mem[222] = 144'h0745fbc4f51108360ade0d5afe580458fa14;
mem[223] = 144'hf063f996f76000ed01ff03b805b7fd6ff136;
mem[224] = 144'h03b8f3d00b4af4ddfcb1038df5d8f05405ca;
mem[225] = 144'hf78f0b5effb7074cfd1f076c00b5fba400e8;
mem[226] = 144'h0504f40afc9a04c1f60f03eb0586034c0bc3;
mem[227] = 144'hfe96fc9bf17905a4f255fcc40d8df39c07d4;
mem[228] = 144'hf225093bf172006efc0d028009220dccfa19;
mem[229] = 144'h05abf66cfd1efb9efee6f1210e2af48505b7;
mem[230] = 144'hf53e0ce10f4df22e007e03e5099cfd80091b;
mem[231] = 144'hfcce02950e9cf07af020f5b1f338f4620fe9;
mem[232] = 144'hf1dbf63bf2cf032bf8e50ca30d63fc21f0cc;
mem[233] = 144'h034c05d209a00d43f1a6f4f3f2b0f2f508eb;
mem[234] = 144'hfcd7f9530561fe4efaacffc6f83902bb04e5;
mem[235] = 144'hf433f2e6fe4605450322f2ea0905f9c10a15;
mem[236] = 144'hfc3afab2f22bf0cd0293017803450909f9c5;
mem[237] = 144'hf96ef733076d0557f880f3cff172f9eb0ffb;
mem[238] = 144'h04ab0844fb4600eaff98070e006af854f37b;
mem[239] = 144'hf267ff2607e9f6d5fa6805ad073bfc31fcd9;
mem[240] = 144'hfcbaf8d90ba30cc1055cf1b1f479fe62fae2;
mem[241] = 144'h0f8cfba1f070f374fc230dcbfd15f04ff7f3;
mem[242] = 144'hf76b0babfdb40989f0ed09be03ccf5e30293;
mem[243] = 144'hf7c5fad1fe240733f425f915f8c604c90bf6;
mem[244] = 144'hf91802d90808fc29f54b0cf0fb2903b30f62;
mem[245] = 144'hf07205bb037c0c310c8cf223f776f371fb6e;
mem[246] = 144'h01f8039c032200d606b60e3afe2903f204da;
mem[247] = 144'h014df339fa950251fdd2f0760c9ff8dafc80;
mem[248] = 144'h0f450515f7d9f98903e5072c08980735feec;
mem[249] = 144'h01530550f029ff4c0d7cf05e0f680e6f05c6;
mem[250] = 144'h09deff4fff0cfb7705a708d9f9650ad4f819;
mem[251] = 144'h070bfa4b05cb02320413f45d0a4df9fcff31;
mem[252] = 144'hf78602fff295fe1ff93702de0a3804c4018d;
mem[253] = 144'hf680ffb9098c01f7fd5e0b72f6810506f188;
mem[254] = 144'hf52cf26104d2f13af734f558f6cbffeb0c03;
mem[255] = 144'hf2e6fd67fd87024409bdf678fbf8011bfb18;
mem[256] = 144'hf6090faafdc80abcf85afdeaf633f59afa29;
mem[257] = 144'h05b6f94efa84f2c902bd0b67f509f4d30f68;
mem[258] = 144'h03e60888fd88f70df413f353f038f2cb0408;
mem[259] = 144'heff5fb42f51f05f10f69fa0bf719f5fc0ed3;
mem[260] = 144'hfdd0fdf50656f00df9cc08ad08f9f8430c59;
mem[261] = 144'h077df3340ee60995f830f0880624f6f6f4cb;
mem[262] = 144'hf4a8f731f042fa740f96f35ef899f107fb46;
mem[263] = 144'h047502df0541f1a3fc15f61900bb07fe0c91;
mem[264] = 144'hf21ef507f4370ed4f77ef8fa0aeff3b10404;
mem[265] = 144'h032b0d2df213fc90f84f01b3fe8d00fb0ae3;
mem[266] = 144'hf0fbf807f5fefa10fcb4fb35f8cafcb50db7;
mem[267] = 144'hfdcbf61800530bb0fc0ef49a010304240f0e;
mem[268] = 144'hfe0cf23e0518f068f1340db1fd53fef8f85e;
mem[269] = 144'hf937fcb30a0202960e52fcdbf752f344f8e0;
mem[270] = 144'hf22809d2fcc1f835feeff0380945f2420dc9;
mem[271] = 144'h0c04fb61040f0f7606d000510c200c06f998;
mem[272] = 144'hf3e9f3910f3701090323f852f3dcf9320d91;
mem[273] = 144'h02480e370504f4a7f9ba0b520550fc31f6c0;
mem[274] = 144'hf22e020ef6f30b72f412072307aef9b9f378;
mem[275] = 144'h03a1fbe80212097ef2e106fbf80c0b3d0f53;
mem[276] = 144'hfe9001970d6606f6f8a20688f17c0431f0ba;
mem[277] = 144'hf186fe0f0b28eff805880360f43bf701f172;
mem[278] = 144'h054f029cf7ebfab7f4c10bc606eefe07fac4;
mem[279] = 144'h05fcff10f09a031c0f84015509f0fd0900c1;
mem[280] = 144'hfc7dfc2506b40d4bf5ab091a0f9903500472;
mem[281] = 144'hff550357fb1600670df9fc83084809d2047a;
mem[282] = 144'h05bdfa36f0eafe50f4180c51f7dd096dfe03;
mem[283] = 144'h00f8fe9b080df943ffb4f9c6f5cff7f8f6e6;
mem[284] = 144'hf0e906c308a505faf47df4970af803d203ad;
mem[285] = 144'h011007e1048ff26406bf0a34f0dcf61efba8;
mem[286] = 144'hfe9208f508affa4a0087f358f55ff7030a8b;
mem[287] = 144'hf260f807fbcbf9170a1d0ebbf492f15d07d1;
mem[288] = 144'h069cfadb0885f900fca100030036fb81fb84;
mem[289] = 144'hf139fc47001cfc4805a007eb0f240af7f7b4;
mem[290] = 144'h0eedfc77ffe50cf3f41b04be0fbcf763f6cc;
mem[291] = 144'h0518f3b10a1500f205f50e3af7e70e140d5e;
mem[292] = 144'h0f56fb4b0d15fb0af9d4fd84fb4a06410ba0;
mem[293] = 144'hf7c6f3eafc2b02cf00e5f88ffe1df6f50a01;
mem[294] = 144'h0ca0f420f9bc0755ff140879fc91fa53f19b;
mem[295] = 144'h04fb0a1d0b7803b3f853f9d407e4f488f288;
mem[296] = 144'h07b3f4cbf04704c808c0f72c07ccf76c0001;
mem[297] = 144'h0fd3f750fcd80d470483f5a007cd013e080b;
mem[298] = 144'hf7fd038f00c70f7a03b40439f9b5f91f007d;
mem[299] = 144'hf3daf68306f1f04afcac0b6af885ffacf68d;
mem[300] = 144'h0a89fc18f63504d4feadf0b9f481effd0f8e;
mem[301] = 144'hff6a029ef32ef86ef409fbc1f8a0f4a8fb66;
mem[302] = 144'hf058f6f9f3560355f390066705d305dd0dd6;
mem[303] = 144'hf093f74c05380b47fa6d0adb0793fb3f0c0b;
mem[304] = 144'h07390551fb33005d078a0fa9f4e6084ef82e;
mem[305] = 144'hf4fb0c560aa8fc51f0540c0d0a2d0118f8d2;
mem[306] = 144'h0384ff82f146f9580dedff30f4180d18f129;
mem[307] = 144'h0504ffe1f2bb08260dbaf2b5f78ff34df8fd;
mem[308] = 144'h0da90fdd09c604fe02a90ea5fb6cfceaf7d6;
mem[309] = 144'h0742009af8bcfcebf15cfef5049cfe280c4b;
mem[310] = 144'h0573f1f6f7360a98ff2d05bdfc6509790b6b;
mem[311] = 144'hf69e0256fab90902f671f6660c6d0773fd53;
mem[312] = 144'h0622f1af03c9f5950acf016af1a408f1fcc0;
mem[313] = 144'hf9e5f49afde70543ff1f0919fefb064d05eb;
mem[314] = 144'hf9ec075afc3906a9097a02b007caf481f357;
mem[315] = 144'hf9fff48504adfd9cefff04ce014afb8df474;
mem[316] = 144'h0c040d6bfd9c0165f57bf51001c50a1c0c47;
mem[317] = 144'hf1d9fdab00aa035a0d120b85fefff844fc26;
mem[318] = 144'h096200cb0e63f38bf6d60d1e0ad0fc970f63;
mem[319] = 144'h0377f2c90072f5cbf910f715018dfcc3fcfc;
mem[320] = 144'h0f070523faee051bfae7f828f528ff2006af;
mem[321] = 144'h00cafc80fb0d0909f475fab30bf309af090f;
mem[322] = 144'hfc440c5b020c0739f8bc0dd8fb850df4fe35;
mem[323] = 144'h059d09e9f742001df488f8ebfd7df963f1d4;
mem[324] = 144'h031efbad0ffdf56a0137082af425f631fde0;
mem[325] = 144'hfdb5f7f60a7cf0fb05aff592f287f9c1f031;
mem[326] = 144'h04a4f63f06f006a3fd8c06f003210b28f236;
mem[327] = 144'h0e4df6810d350134f2d4ffbe09c90530f05e;
mem[328] = 144'hf01405e20ef7f5a904fbfa7af067f9a501fb;
mem[329] = 144'hf870f54cf5c3f2fa0905f9adfe1a0f54f066;
mem[330] = 144'hff760fb401aa0fd502d20770f71f07860661;
mem[331] = 144'h005f0985f297f74d07b408200493f10502c3;
mem[332] = 144'h0e1e03d704b40662fa4e0cf00e8502570bf1;
mem[333] = 144'hff2d0e64f8d0fd31f5e7f8f8f52a0a580637;
mem[334] = 144'h042af9ecf66cfab40551f5510ca00293f98e;
mem[335] = 144'h04bbf64004f2ffe80e0af34ffb3ffb3efacd;
mem[336] = 144'hfe330c2400aef84bf66c0966fa3cfe9503dc;
mem[337] = 144'h0cbbfadef804f378fab90b7bf459f56efce8;
mem[338] = 144'hf0f90cf6f192fadc0e2af316f61df105fa73;
mem[339] = 144'h0b2dfae7f7dd0d060c4d03130a68097c0a45;
mem[340] = 144'h02ad0eea099f03e0094dfbb60f6ef9d3f455;
mem[341] = 144'hf006f4faffbbfdd6f98b09e600450a0ff7fd;
mem[342] = 144'hfd14f72e04bff50fff980359f0740d6405e5;
mem[343] = 144'hff2dfdcbf7d1ff1bf4620363f6fc04320cc7;
mem[344] = 144'h0148f21502b9fa61f715056f09c2f93f0269;
mem[345] = 144'hf67607f4f1a50dabf03100bd0997f2c4f78a;
mem[346] = 144'h0a78f0a20e2ef4460212fb2b0055f1f20369;
mem[347] = 144'h00b9fecb02c8fe4afbd6f3ee029cfcb4f8e9;
mem[348] = 144'hfcbb004f0e61f753f5d40f850bf90ea60821;
mem[349] = 144'hfb44f14306de0180f952fbb40ee2f3b30765;
mem[350] = 144'hf74b01320f1b04720b6ffdf6f288fcff0b10;
mem[351] = 144'hf160f0f20a36041efdbb0572f86efd2cf97c;
mem[352] = 144'h0dc2f85b0691027afdaffceffb51f874f926;
mem[353] = 144'hf3eff342fc3d02abf192f7d80b9e06cc005e;
mem[354] = 144'h0b71fff20be9f8b9046b032b06dc02fff931;
mem[355] = 144'hf12dfff4fb43f3f4f0a10a8203bffe22f5ab;
mem[356] = 144'hf39ef0cafa55fd96fbed019efd4d062cf6e6;
mem[357] = 144'hf705fd7eff01fd2df34df093f7f302aef193;
mem[358] = 144'h04fb04800da90f3e0fbbf451061af95e022d;
mem[359] = 144'hfec4fdd9f27cfa9d0dbb09d8f4da015efbfb;
mem[360] = 144'hfcc60245002704440273065805ee0c4c07fd;
mem[361] = 144'h0b89f26a0db8f73af4b2f9e7032d0e5bfa83;
mem[362] = 144'hfdc30ce501e1f087f5c90ae503af066400c7;
mem[363] = 144'h01ef0ea3f91f010f0618088405d003ab01e9;
mem[364] = 144'hfb6d05c506e2f4e70a76f7fcf9360e930612;
mem[365] = 144'hf401f6c5f744087903ea0c19fa19f80bfcc7;
mem[366] = 144'hfae0062f001ef4fef255f95a0476f66103a3;
mem[367] = 144'hf5daf19407cdf2cafaa007370bf2038306d9;
mem[368] = 144'h005b08bc08b5fa72f95d077b0d4bf55c07a1;
mem[369] = 144'hfa6c0a03fc80f59b052d0be8047a05cd0035;
mem[370] = 144'h035000ef0b85f5720bebf779f5b1f166ffe2;
mem[371] = 144'h05c0f3c5fd160b45faf708fbf634ffc1f119;
mem[372] = 144'hfcc608e4f0cd05aa0810f715fd01042b08ca;
mem[373] = 144'hfc6b01e0f49a0c51fee90069fc020bdffb1d;
mem[374] = 144'hfcbdf706016001e9f28b0227fed90cdcfda5;
mem[375] = 144'hff590be1f911f8f909e003af086bf80ff061;
mem[376] = 144'hf9df0e64f4ecf90c0ea3025b0d8dfa7ff3cd;
mem[377] = 144'hf41bf25e03430a7f05f00c0afda9f18dfb3a;
mem[378] = 144'hfa15077af34607b6005ef22bf85b033304e4;
mem[379] = 144'hf9a50d06f94402e2f4e800e309cd04fd0417;
mem[380] = 144'h0c01f287fb3ef4fb0b3f0e91fbad065d05ba;
mem[381] = 144'h0746fe2af45cf6ccf1fffd95fdfb07c405c5;
mem[382] = 144'hf8a1f1870038f777ff5bf3ebfee1f8ebfff2;
mem[383] = 144'h07760a5d07770bb1f77f050806cc08b2f808;
mem[384] = 144'h03800bbd0f0bfc5bfe33fabc0aae099d06fa;
mem[385] = 144'hf2b2f46af78df5b5018efc22056bf81af21d;
mem[386] = 144'h0b1e0d19fad3053ffbbff1040f94fd98f5d0;
mem[387] = 144'h0220026bf399f599f7a001c209dbf0f10882;
mem[388] = 144'h0e2cfe150773f5b804e1f830090bf7fef2ca;
mem[389] = 144'h0733f9a9f313f713059e0d2e02d00778fbcc;
mem[390] = 144'h030c059cfdf7ff0bf03cfaf108b7f2fdff5b;
mem[391] = 144'hf4cb07e7f9b10b360bb9fcee0ef9f2560005;
mem[392] = 144'hffa4f38a052bf9a4fa2506370af2f419055b;
mem[393] = 144'h0a35f82d0e600d8a012cf2a1f9fe0e61f0d0;
mem[394] = 144'h0661f533f723f6120ed6f4950d23f1130fa8;
mem[395] = 144'hff82fa9bfea90666f3630b47032ef69900b5;
mem[396] = 144'h0feaf211fd700137fbb706faff48091e007b;
mem[397] = 144'hf60a066ef81d035c0aa2f20c071b0fc80f58;
mem[398] = 144'hf86a0eb50b460be80847f485f90408310c27;
mem[399] = 144'hfb810b9105990a4004ef0e90f80cfc7dfe20;
mem[400] = 144'h04d0fe84f00e000efac5f009f272095df196;
mem[401] = 144'hfb19f9280f77f9dc0e630ccf09de073a0835;
mem[402] = 144'h0020027c0f1f0125f78e028ef08600a70dd8;
mem[403] = 144'h0606004efcd108740f81f11d0f50024a0143;
mem[404] = 144'hf6db042dff210c6201960779fddcf163fccf;
mem[405] = 144'h0853074ff9860f1f08e107d80fb406660659;
mem[406] = 144'h09a004f4043bfc930f6d056dfa6bfc9105a1;
mem[407] = 144'hf3a1fc7703aef6a80b72fee90cd6fc4cfe17;
mem[408] = 144'h0fc701da06750c76f40d0cbe026000d60b0f;
mem[409] = 144'h0b40f4d3013209dd0167ff3af9d1f61efc51;
mem[410] = 144'h01360e1d0856fb5a0179fca5f2660dc9096b;
mem[411] = 144'h09a0fed1f198f08df19004dc0f82091c0bae;
mem[412] = 144'hf544f4a1f574f26cf3860da5fafe008afd90;
mem[413] = 144'h01a0fe02f6da01a00c3f0dc9050cf49ff942;
mem[414] = 144'hfe910ed4f12cfbeafe60ff8bf21dfec209a4;
mem[415] = 144'hf88dfe68f09df1b609f8f060fe61001a04cc;
mem[416] = 144'hf52e0a5d0a82f06800d4f6e00ab8f75afde9;
mem[417] = 144'hf33df20206950d14f3fefbef0a43f5180176;
mem[418] = 144'hf04008d30e8d0a88f5fe0af3f1460ae40e15;
mem[419] = 144'h0ca8fb5e05a1feb20b17056bf4c10251fa9b;
mem[420] = 144'hf574fa0cfc90f51e0b3afa180270010102e2;
mem[421] = 144'hf7b3fae20f7800500a7b08f2f13a0b56fe20;
mem[422] = 144'h05d1f9b5f70bf2b30e67fadaf52f05b2f680;
mem[423] = 144'h05dff553029df453f72df03bf63a0e8c0b47;
mem[424] = 144'h0e93f43a02a40f5207afffac0895f6d2f907;
mem[425] = 144'hffeaf6180ef10721ff72f3c10701f673f619;
mem[426] = 144'hf434f79ef1c3f90701bdf22cffd40f32049e;
mem[427] = 144'h004d0d12f215f34d00f9fdb3f65ef8ce01a7;
mem[428] = 144'h0d390284fa140dd8fdb4f7a5fc270dee06ee;
mem[429] = 144'hf6e00150013b04b70e50f5f3f8b605330e80;
mem[430] = 144'hf683f402f8b3f76bffc9f041fb75044709c8;
mem[431] = 144'h07cef7070c530b40fc03fc7df127f136fe8c;
mem[432] = 144'h0426f65c0748fe200f3d069cf977fd9b0b6e;
mem[433] = 144'h03f50f80f9bff542f28bf27af846f8180ded;
mem[434] = 144'h0d6805280fa2f88e017301cb09bd03f902ed;
mem[435] = 144'hf87d0b7701550364096c0b2a0b3a0797027e;
mem[436] = 144'hfb190d7f0b85f321fd9afd8404d0f5a3f649;
mem[437] = 144'hf105f133f25a0a36fd8afb81f84ff4140c1d;
mem[438] = 144'h0ec801e2f177f8c008e9fa54027cf4b0fbc0;
mem[439] = 144'h0b33012d060201da05d5fdcef4abf094ffdf;
mem[440] = 144'h09f3f35703130b260d81f8460b460cc40866;
mem[441] = 144'h0bc5047ef507f463f350069005cbfaa9fd60;
mem[442] = 144'h08310df104bdfd1ff62e088df0e4004f0c49;
mem[443] = 144'h0a38f64a0f1a045ef47e08ef0b5dffe00f73;
mem[444] = 144'h0f8dffe3f4b2f4b60d600457f9b705effad4;
mem[445] = 144'h09d5fef60477fde0fb240f410026f3effeac;
mem[446] = 144'h0fb2fb7605300a4206efff170ed2f7c6f252;
mem[447] = 144'h053ff24e00aa0b6b0e480e05f6590294f5eb;
mem[448] = 144'h0c2a0a250d20f082f3060c30f2640dfd06d3;
mem[449] = 144'h0f61f144f5f6f121fba7f73604d7faea0694;
mem[450] = 144'hfd24ff07f50bf5a3f8290ae00b82f827f006;
mem[451] = 144'hf21dfae3fb60fba60ccff217f79bf2690b58;
mem[452] = 144'h03d8f725f1d6085d026107f3f10e00b3064c;
mem[453] = 144'h0e3dfcd3f82ff67100000e99f96ff3edf682;
mem[454] = 144'hf90b04adf683fba8f240f6a6f7a8f1e00850;
mem[455] = 144'hf467f069f45c05c0f95ef4e5fec102b0f35e;
mem[456] = 144'h0eb40979f086ffc7fba705cffc63fd4bff3b;
mem[457] = 144'h068108fdefcc070001e701440178f085f9b0;
mem[458] = 144'hfd26fae3f5630a22f89efcde0112f494f6e2;
mem[459] = 144'hf29105fa0c010ba8fb76f71dfd3df4740842;
mem[460] = 144'h094cf4faf57effce0003039bf21006fdf338;
mem[461] = 144'h0c460a4d01f008ddfde4f4e20f25f7abfe5e;
mem[462] = 144'hfabbfb5b0e600b5c0510fde7fe1604a903fb;
mem[463] = 144'hf90efdb5f9c7031105500a1f018df6eb03b2;
mem[464] = 144'h0de8f013ff40f345f1d40eb1f94406e4f63c;
mem[465] = 144'h04b7f6d4fca1020b01f60be50b7e0e73f1ae;
mem[466] = 144'h0767f6f0f017fdccf9c9f68a021a0cf30ce4;
mem[467] = 144'hf9dbfe8f0512fcdc08f6fb8bfd5309280460;
mem[468] = 144'hfdf1fbfbfc4e0c9c0895fb4cfced0be102f9;
mem[469] = 144'h00d6fa3ffb6ef6140426fb31f675fe72f32e;
mem[470] = 144'hf05505400b6c0976fd3bfbb8f30df339f321;
mem[471] = 144'hfe22f3ccfb1afb880870fed60cf10c220922;
mem[472] = 144'hfab40c8b07d90bfdf3c40aa3f3abff66f522;
mem[473] = 144'h0409f02c0b610897faff0e370bfffb7f0434;
mem[474] = 144'h0830f7ac0072f6a90db8ffadfbb8f536fd90;
mem[475] = 144'hf727f9e10ac1f7550b0107effc56ff140733;
mem[476] = 144'h0a2cf597faee0bc3f44302c2fe0bf6450fc4;
mem[477] = 144'h024c0c1f0e90f39a08b10b75f5b80ddcf776;
mem[478] = 144'h0be607f20f12f19df7c60a8204a9fee2f2d1;
mem[479] = 144'hf87e0752f512ffb7fa2709a2f128f9b5fee7;
mem[480] = 144'hf75f05b3049b0393fab8f08603b6f2f90fa7;
mem[481] = 144'h0720ff4c0920f2e7f5d8f6490258fc24078d;
mem[482] = 144'hf4ca0326f7eeff37f07a03d5081d088405d6;
mem[483] = 144'h0914f79605a4075c0ac3f828fa4ef62bfd55;
mem[484] = 144'hfd4ef9dcf489f7ed0142fe490eaf03a2feda;
mem[485] = 144'hf4eafb6904740c42070a0bd10436f93bf754;
mem[486] = 144'hfcecffe6f375f02cfb3efdf2fd0df3000439;
mem[487] = 144'hf074043803e705d10a5509e7f5dd026d0dbc;
mem[488] = 144'h0bfef92b05520690f4f20efbfe1af26c0852;
mem[489] = 144'h04050f56fa1e05c60a2f0586f205ff88f553;
mem[490] = 144'hf50d03a1f8f5f439f32dfdc0f597f3870f05;
mem[491] = 144'h087906f30cb4fd9cf442fdc6fe0c0ef40d6f;
mem[492] = 144'h01e9f56e0743f9f9fea00c2c01d7fdc5067a;
mem[493] = 144'hfdbdf0ab0862fa3007b10476f46ff43808dd;
mem[494] = 144'h0e4f0ae103b8ffb00c400187fb1cfea1f55f;
mem[495] = 144'h0656f080f40302aff11c0a6d0be40fb2fb18;
mem[496] = 144'h03800a52fbe0f5b5fab109b0f3f20dce040c;
mem[497] = 144'hf94dfc9df738f6b3fd880d9504200b63f0ee;
mem[498] = 144'h0a15f5e5fb14092002ccf591009e0200f25c;
mem[499] = 144'hffda08a2f4340e90fa46fdd1fdde00f30178;
mem[500] = 144'hf920f135f176031c0f7ff115030ef8aff7b7;
mem[501] = 144'hfb86f1a3f30f0757fd0f075b06db05630389;
mem[502] = 144'h0b4ef0eb0edaf7460f69feda0a44fc970828;
mem[503] = 144'hf2d2ff7c0b6efaeb09370158053c06d70b56;
mem[504] = 144'hfbd9020cf0410e6c0ba00bd2f6eb0eba0ebb;
mem[505] = 144'h0d67f026f6350e2bff19f8b90c77f598f34d;
mem[506] = 144'h053b0d9904c90ac8f5db05c3f7c4fe7a050f;
mem[507] = 144'hf1bdfbe6fbec0f7cf6880869050bf8350be9;
mem[508] = 144'h0558fc0af9faf1240d88032c09b40fac009a;
mem[509] = 144'h0465f925f1f20edb0845f9bc0ca9f2df0adc;
mem[510] = 144'hf40af8aa0879069b0ab1043900d6fd0af927;
mem[511] = 144'hf5dc014afc9bf28e0842f25d00eb0db60680;
mem[512] = 144'h0efa06cdfd8906d7ffd4f3e70b83fc1a0bc6;
mem[513] = 144'hff59fe400584fea3f693fd14f9970286f888;
mem[514] = 144'h0d13f63cf773f42d0ec9f93e02b90cb10fdf;
mem[515] = 144'hfde5f888fe0b0c1f07c2f9c2fa660d5bf5ce;
mem[516] = 144'h0cf6035d0655f272f35d07450ddb0b58fd35;
mem[517] = 144'hf8b507b5f0c007dffb4bfd6e00fdf72f0304;
mem[518] = 144'h0ef6082afcdb05c30dd4f858f4fd0f4a04a0;
mem[519] = 144'h05870fa5fefd0a530359f134fe4106c5f4c8;
mem[520] = 144'hf59af06704b5f80eff72fc50f3abff25f778;
mem[521] = 144'h0f4b09c50fd306af0f3ffebf03d00a5ff98f;
mem[522] = 144'hf3220452fc5d05bef7bcf4c2021f011c031c;
mem[523] = 144'h05c2075706d8f575f6c6f4dcfffefe84f6d4;
mem[524] = 144'h037af9b100fdf7d70136011e005cfb9ef2ba;
mem[525] = 144'hfb2ef253034e0b60017ff09bf654f2f9fe8b;
mem[526] = 144'hfd440cacf9a202000eb60aa5fe2e080f01e1;
mem[527] = 144'h0029f0a2f1d5fa870e580ae70f70f889f32b;
mem[528] = 144'h0a35fc6809fe0e2efe08fbb1fe43f5fdf4bc;
mem[529] = 144'heff9effffc89f683fc79f3aefc1c00dc06eb;
mem[530] = 144'h08e20b93082ef1a40b31f096f619fbc4fa0d;
mem[531] = 144'hf56200c90dea038205430eedf3290f8af788;
mem[532] = 144'h05d90abf0d3bf887f9a103e20dfcf50908a7;
mem[533] = 144'h0273f27df9dbfce7fa45006ff25cf6ac0107;
mem[534] = 144'h0a00090df5b4f126f0740c73f68c0227053d;
mem[535] = 144'h0e090501060d051df48ef8e30984fc09f288;
mem[536] = 144'hf7ecf99ff47d0d8bf665f229f21cf56af187;
mem[537] = 144'h054ff366f6a9f7d3f1fb052df1e9f0c1fa12;
mem[538] = 144'h08a80f50fd25f7d007d103b5f2150a37f9ef;
mem[539] = 144'h0be1f1ff0f6306e2f7defab4f08005130562;
mem[540] = 144'h0a9ffddaf8a5fc280b230bcaf62efa6b0d15;
mem[541] = 144'h0da10f69f5dd0bda090d0e4ef2520962fd68;
mem[542] = 144'hf6dff111fccc0b1ef5aaf7d405c0f321f7c4;
mem[543] = 144'h063cf5b3fb760ca3011cf65efffff4adf60d;
mem[544] = 144'h08d1f055f47d07070c2b07bf08290289063a;
mem[545] = 144'hff5c052304bcf499feb4fed4ffeb0fb4f475;
mem[546] = 144'h083af405f73a0414f0400671001cface09e5;
mem[547] = 144'hf87500d102260ef7f940f42805770f0ef689;
mem[548] = 144'hf35602d2fc460b15fc27f405082ff84df121;
mem[549] = 144'h0479f9260e590718fecbfaa7f4bb034a04b1;
mem[550] = 144'hf5e80a2201dc0929ff1ef183f2e4f8cc02c8;
mem[551] = 144'hfea60ef9f2dafb2c0d51f1870354f4bd03ed;
mem[552] = 144'h02680cec04bd0820f7fe02afffbff1acf364;
mem[553] = 144'hf49a0d3af88cf5bcf6db03b10f350522f0f0;
mem[554] = 144'hf09e09a9f221048ef7ce04b3f6740afdf043;
mem[555] = 144'hfb940503f01cf0d1020506ef04b5fd3bf20a;
mem[556] = 144'h0cd50c4400ac0d15f852fd9dfd640c01fee8;
mem[557] = 144'hf7a5fabfffd0f8b50adf020f08f0f43e0480;
mem[558] = 144'hf9f6feb600e9f399f1e4f89f0f7f0c1f09f0;
mem[559] = 144'h0c4cf057fd4bf1550e71f3eef16ef49ef55d;
mem[560] = 144'hfbd3f67ef7c9f706fad9f3ef04b103f802d9;
mem[561] = 144'h0d2cfb00f1f7f62e0f6c07fef6bbfc830f30;
mem[562] = 144'hfcf704a8fe59f0ee04490e77f1a103cdfec4;
mem[563] = 144'h05e20bf2027c044afacbf6f5f194f9c0f84f;
mem[564] = 144'hf2abfba1f7c705e3ff20f6e5013e05750371;
mem[565] = 144'hf3cdfd540cf8fd56053ff3aa05e003980847;
mem[566] = 144'hf145fc40fd3205260cbdfe5f08a4056507b0;
mem[567] = 144'h0ead0c2ef1d7f29cfd8afb40fd8ff50af31a;
mem[568] = 144'hff0202fefa9e05160680054ffc2509d309aa;
mem[569] = 144'hf111f0ef0e59f859023df3170ca40749f858;
mem[570] = 144'hf934ff70fc25f1fdfd2a0da90ad9f9ae0f84;
mem[571] = 144'hf0f7fe73fe79f5070b10fc42feb5fa84f2f3;
mem[572] = 144'h0a08fbdf0f160b4ef215f0b5ff320b21018f;
mem[573] = 144'h0e92f4e9f802012f009af83f0c00f34806e2;
mem[574] = 144'hf03302fe0dde0999025c0a290ee508dff23c;
mem[575] = 144'hf049fde6f63ef8690450f8e90896f4440c5e;
mem[576] = 144'hf04af4bd0ee3f3b7f934ffdbf6c2fdc8f4ef;
mem[577] = 144'h073af665fcc7f008f24e03d8fb4606f00759;
mem[578] = 144'h0675fdfef84df45bfb7f07f7f1cbf2c702c9;
mem[579] = 144'h09eb0dd3087708df0d130c6df649080e0e2a;
mem[580] = 144'hf06df4790d06ff98f71ff9de0a60f73bf28b;
mem[581] = 144'hf0c60635074a0f92048408fdfa7f0fabf9c7;
mem[582] = 144'h0329fb2309340829f4730c6e0f4c03a8fed7;
mem[583] = 144'hffbc06530a360304f3eaf44bfe9efea0f0e1;
mem[584] = 144'h072b026c04a5f719085bf864f51cf044fc76;
mem[585] = 144'hf6a10340f050f250f93a0783f980f1a3fa71;
mem[586] = 144'h069602c500e506d5f878f21b072a0bc3f6fd;
mem[587] = 144'hfab2009bf93c04e10198f250f8680aa20db6;
mem[588] = 144'h0babf242f1f2070b033dfd39face034cf11f;
mem[589] = 144'hfdf506a8fdd600b6ff12f5200117ff420a0f;
mem[590] = 144'h02bc04bef655fbd4fdb7f534f9abfbe90cbe;
mem[591] = 144'hfc05f1e9f95706280295f968f812f2a1f35e;
mem[592] = 144'h04af0363f949f8c5095ff6d2f9d308a00125;
mem[593] = 144'h014a0ad80c5904c807f103e00582f2820793;
mem[594] = 144'h0212036cfb100639f3a30837fab6fc04ff47;
mem[595] = 144'h0686f174f7e70cc0f10803dbfff3f69a0479;
mem[596] = 144'h0d66f3ba0676fb6afa3ff0fdf0580a6efd4a;
mem[597] = 144'hff48f75704f9013ffb00ff360af10f9df956;
mem[598] = 144'h0753facaf2620091f7e00d28fe340d4ff46e;
mem[599] = 144'h08f5f292f2e50cb3f258fb830e04f11cfa44;
mem[600] = 144'h0a3b0bb203870a3aff8c044c09b9f64f0218;
mem[601] = 144'hfab0071c0c4af0fefb320b57015e03600eec;
mem[602] = 144'h09f809b0fe6e0febff0c0e5308430033076f;
mem[603] = 144'h01620a4803970371f7e1f1850ec000d403aa;
mem[604] = 144'h0ea30599f7fef3c7fa2a01bcfe7cfea4f3c6;
mem[605] = 144'h0068f8fb0001f701fe19fe230190f293f0d2;
mem[606] = 144'h0049047003b90fa8f21e0f10f64afbcd0762;
mem[607] = 144'hf9fa0689059efa46016c0c4cf76c071100b0;
mem[608] = 144'hf9720d5df5af00910a6d0725fe54f3b2f62e;
mem[609] = 144'h0d850d390bdb0843facc0c470d84f24e0135;
mem[610] = 144'h028a07980ce3007f01220121042ff5ee01a3;
mem[611] = 144'h026f0f4005f8f7400645fcbcf8cf0b540a56;
mem[612] = 144'hfbc30f660ca9f6d3f742f67107e3fa5e0f89;
mem[613] = 144'hf4ed0955037cfd5302a0f45b0e1b06e5005c;
mem[614] = 144'hf195061af0a10f74f3f4f4ecf3f4f65ff9f8;
mem[615] = 144'h055dfe1ff66b0e420201f63b0cf707030469;
mem[616] = 144'h09540a7a09aafda10d50088eefc70681f475;
mem[617] = 144'h01c6f23f04b3ff40ffd5056efaeaf00dfda0;
mem[618] = 144'h06d7fc4102e106c7fc14f162fa4f0235099d;
mem[619] = 144'hfda10f31fdf504dbf647f727f0020ec50666;
mem[620] = 144'hfc590e82f6b5feb8f7420730f277f63bfe38;
mem[621] = 144'h080602c0f18efb8e0699f587063502bafffa;
mem[622] = 144'h0323ff5706990bcc04cbf82f0afefda6f637;
mem[623] = 144'h09310315050a02c8f4800361f3430b7dffc4;
mem[624] = 144'hf79b04d0f08f0e47f515061d076b0e3407b3;
mem[625] = 144'h0ea60012fccefaed0a990e5a0e43fcac0923;
mem[626] = 144'hfafff9b4f068015cfd32f8d30c8909eff59c;
mem[627] = 144'h0fc30433f943f33df6aefb65fd6a04dbfc57;
mem[628] = 144'hfd8101550e55f752f0b2f228f34cffa00af6;
mem[629] = 144'h0dae084df6a7f23e0af3ff6507e10a5206ec;
mem[630] = 144'h09a3fc4b0ad3f5b0067a02aaf7c5f1760b12;
mem[631] = 144'hfbfff004095cfdc4f460f94e035c07fc02ad;
mem[632] = 144'hfb72f4aa0c3ffc6b03b90487003fffe10026;
mem[633] = 144'hfcc8071a0e77fcef0ca7067bfb8004b60750;
mem[634] = 144'h0a2e05110ef20eb8f6aef5650703f4480337;
mem[635] = 144'h0804ffcc0c23fe4d029f0886f4d10f1d0ec0;
mem[636] = 144'h0374ffa3f8d7fc9afc8b04b6097c0d8af598;
mem[637] = 144'hf646f7b1f5bc04c307eaf2260b77f4a00c29;
mem[638] = 144'h0c240202f1780b790674f3350167086e055e;
mem[639] = 144'hf3b8098407710901fd660cb4fd7d020a0ac9;
mem[640] = 144'h0e40f82f0837f550f07affbf0c00f2c5f950;
mem[641] = 144'hf1280080fb61fce6fc790898fd61fb9f0d12;
mem[642] = 144'h0678f15ef43609de0058f7a1058a070602c0;
mem[643] = 144'hfeaef24a02070a810a5c04ae0305f309f55d;
mem[644] = 144'h026cf2c40df90879f07df000f18c0870f1ad;
mem[645] = 144'hfd04faab06680af4f5800cc9f0a1fb9b0d1e;
mem[646] = 144'hfc80f095f3aefdddfa71fe190b7406490508;
mem[647] = 144'hf223059105940d46f3b407c80be4fe33055f;
mem[648] = 144'hf494f18106f1ff11f6fa046ff8c30a270e3a;
mem[649] = 144'hf1570d13fc23fecaff7df2d90034fe00f5f6;
mem[650] = 144'h0c360383f2fd091cf26f00c8f6c50d93f4bf;
mem[651] = 144'hf8bf03a3fbd7f61e00f108fe00e8f37a09ba;
mem[652] = 144'hf693f40a0a32033c0520f935f69af04ffc55;
mem[653] = 144'h0c250db8fe0ef8c709a3fbd20ba30cecfe92;
mem[654] = 144'h0428091702be0f3a034ffe660bea08c100ff;
mem[655] = 144'hf452fa23025a0add046704a2fbcafd7700cb;
mem[656] = 144'h0c3e0c0ef8570f28fe93ff78f397f5920ea8;
mem[657] = 144'h078f02c80872fa32f392054a0fc508c90f03;
mem[658] = 144'hf51c0aacfc6709650c5bf92805ed0596f4f4;
mem[659] = 144'hff9df6930420fd95f6fb0766f17502710794;
mem[660] = 144'hf5f3f8310fe5fcad0915045af5f1079b0747;
mem[661] = 144'hfcc8f72ff5cb04d1f948fde407a3f477fa2b;
mem[662] = 144'hf1bbfe610e4303f8f3160ef8f1e9f4e7fc39;
mem[663] = 144'h047c0894fed501b8fbf10912fa26f8fb0928;
mem[664] = 144'hf4c40bdb018cf8720a10f917f99cf5250c9e;
mem[665] = 144'hffd80620030003e6f191fc30097a0352f75b;
mem[666] = 144'hfadb015af1ccf7f80e07f482f96bf034f548;
mem[667] = 144'h0e77fc5806bdf672f452049e0b05042d05a8;
mem[668] = 144'h026a08d8fa8a0e03f150f817f4def5c3f672;
mem[669] = 144'hfccaf48ffb4f08600d8efe3bf7b5faf80f2a;
mem[670] = 144'h0d290a990341f2b602f9f8dc0f53fea4f47f;
mem[671] = 144'h0c890d4e026df9d6f31af97c017c096ef703;
mem[672] = 144'h060e0570ff92f6d60c7c0169096bfc7409fc;
mem[673] = 144'h0a43fcfa08aafedcf0680eba0bea0b7603d6;
mem[674] = 144'hf00cfbd10ae6000ff4c70ed106430d3ffe41;
mem[675] = 144'hf8c4fb84fcc30744f330076a0c5f0ed40bed;
mem[676] = 144'hf0b6f6b6fcb30a53f09809b0ff21045af3ad;
mem[677] = 144'hf4e606ae0c9afbc0f177050afac6090af733;
mem[678] = 144'h03ddf8f00395058ef71508def1ee05790d58;
mem[679] = 144'hfe300d2e0cba0def0fd80fd008b4f48dfc2a;
mem[680] = 144'hfb90fd6f063b02d7f56e093b04d80b09fd59;
mem[681] = 144'hfe390c63f818f95df5a6f1bcff40f4e502c4;
mem[682] = 144'hff21f67b0bc2f03800b4f82dfa1df668fb35;
mem[683] = 144'h0d3dfddaff23fb25f17a07f0f5690af1fb33;
mem[684] = 144'hf5dffb1ff717020700af0520fba60faafb3b;
mem[685] = 144'hf1f2ffe306e3f49bfec7fad6f736f9890720;
mem[686] = 144'hf967071cf5d3fdb006e8fd50f11d060ffdb2;
mem[687] = 144'h05acf71603be0daffd05fdddf44205c4f0cf;
mem[688] = 144'hf060fd050ea60362f9d7f1b1f20a050ef726;
mem[689] = 144'hf3ca0a450122f416fab6f3400009f6aa05cf;
mem[690] = 144'h01f60518f6d0f8d9fde3f75a09940a400131;
mem[691] = 144'h04bafd85f7c60df903d10e7b0b6a0ae5fb3e;
mem[692] = 144'h050efa11051e00cc0ce2fc9cf04df7f8ff88;
mem[693] = 144'h0bc0fcc9f1a00628095cfe7f097d0475f37c;
mem[694] = 144'hf4f2fa68f8330d230af30e5cf82bf1ee00a7;
mem[695] = 144'hf490fb1afcd7efc8fafc0bd0fb04ff8ff24d;
mem[696] = 144'hff86f476015c0ecf0d3af90dfe5ff952fe51;
mem[697] = 144'hf99d030702fbf323fcdb09070f7bf46e0436;
mem[698] = 144'h056b00ed063e015ff8d50c78f62bf585067c;
mem[699] = 144'h0e23fa14f87f064cff430650f27b09c508f3;
mem[700] = 144'h0612fbeff5310368f10eefe701b2092c0b79;
mem[701] = 144'h02b208130a55023b0ef8fd54f38efe470649;
mem[702] = 144'h0511f6e5ff56006bfa0df03dfbe20d810d98;
mem[703] = 144'hfb55f513f85602b3099b027cf6b1f69900d7;
mem[704] = 144'hff4202d8011cf4b40fb90adffc4b01dcf67c;
mem[705] = 144'h0374057cf21bf5b801540680030dfceafa1d;
mem[706] = 144'h01770ca80de8f3d3f1e1012c0522017dfebf;
mem[707] = 144'hfcf508140dcff97df352f177f2a007f4f5b2;
mem[708] = 144'hfead0ceb0a55f349f64af8680b76077f0bcb;
mem[709] = 144'h0bda0dfffa27f8bb0947f379f51c0f87fa4f;
mem[710] = 144'hfa38f152061b0cff090af754fe03f0b7f504;
mem[711] = 144'hf21b013004dbfd9f0cd1f661f9bcfb75fdae;
mem[712] = 144'hff9df6fafce60c16089f0e7a03b10272fa2d;
mem[713] = 144'h0b470f04f64c00d50495f5b6fbb60f05fd7c;
mem[714] = 144'hf36302890b100feafd4d06e8f8920f14f01a;
mem[715] = 144'h03f704fc05b0f30c059afacaf6a9ff14013c;
mem[716] = 144'h0745f579f9d305bdf152f495f9b2f67d05fc;
mem[717] = 144'hf9530e370aa90e040217f4faf4e605ccfbcc;
mem[718] = 144'h0365f249f7de0287fa15ff9dffa8fd1af5d2;
mem[719] = 144'h090ffc6a03f000c305c40c940d10fb780430;
mem[720] = 144'hfc5dfa0df37a0b1cf4e1fb1efa51fd640e0e;
mem[721] = 144'hf36d0bf9f7e70d45083cf9faf08e00effe66;
mem[722] = 144'h01a0f8bc0f080c5ffc31f68d00a2f07f0ab1;
mem[723] = 144'hf9750d3ffe5df9fd0991fd85f5a606780fd8;
mem[724] = 144'hf66600a903eaf18c037df915ff26faddf088;
mem[725] = 144'hf2fa04f20b50f4a3fca5fb27045a08b4f142;
mem[726] = 144'hf8b5019b00e1f20af5f1f20905ac0af10613;
mem[727] = 144'h088d04e60eab035dff05f6be09ed08ff0920;
mem[728] = 144'hfdbcf9eaf54f0ed10d6cfd78fc800f20f311;
mem[729] = 144'h014e09e805de0d44ffa3faf40b1307530487;
mem[730] = 144'hf460f74a032f03e3f877fcc1f1fc03acf4e2;
mem[731] = 144'hf6880520fa7c025ef24c09e8f681f792f7a0;
mem[732] = 144'h01fcf430fb6bf80800390745fef20b1306c0;
mem[733] = 144'h03b9f7d00878f266fb33f4e60cd6f12008a4;
mem[734] = 144'hfcba04ddf257f8fbf7330d460a500817f6a4;
mem[735] = 144'hf785fece04e8f6ff0a94f45e08a60aa7ff5f;
mem[736] = 144'hfab801940635fa56f68ef9b7074df294f1a0;
mem[737] = 144'h05780dac052a0c0107b504670ba4f2e60986;
mem[738] = 144'h06390feafc020f0c071dfde3fa9df3070fe0;
mem[739] = 144'h035f040400ea01970ce4f049f06df7ca0ea5;
mem[740] = 144'hf649f531066a0e0b00bb06d6f4ccf9b00a34;
mem[741] = 144'hfa7ff315f3aff9bcfa17f952f45e0edcfa6a;
mem[742] = 144'h011bfbf503f10463fc74f71ff82407e808e9;
mem[743] = 144'hf57af579f9830919f8420df40091f43cf98e;
mem[744] = 144'hf2910837f72c0067f6fbfe17f8ad0b46fda8;
mem[745] = 144'hfb1f0ebff4a6035a0dc3f25cf0dcf0720c3d;
mem[746] = 144'h0ab90ff30938f87d00c9f14bfd75ff870e7d;
mem[747] = 144'h0b45006a0b9f0a8c0e42f781fc7cf37bf1cc;
mem[748] = 144'hf21afe8ffa5d0129068502f500b20dbaf0f9;
mem[749] = 144'h065505c60b510199f4010cf2f64b054ef305;
mem[750] = 144'hf501063402b7f85c0d32efde0206f0810273;
mem[751] = 144'hfbd400540b22f7f5f06908defdfa0cea03ae;
mem[752] = 144'hf14c0e40fa3803160dcb0f47f34506e10a09;
mem[753] = 144'h00bd0a34ff1d03b7fd3ef6bff4ce0b91090d;
mem[754] = 144'h0dae0ab30f830e29f30bf48d0de400780f1c;
mem[755] = 144'h09510e95045001aefa00068502e1f147f4fd;
mem[756] = 144'h0631f498ffaa03ab069df636f7daf4110915;
mem[757] = 144'h063108fb0800f3940fbdf0290a3ef4aaf37a;
mem[758] = 144'h0b4e0fef03dcff65f84e09010645f31d0b16;
mem[759] = 144'hf6e30f8307320f25f8230557fba207e2077d;
mem[760] = 144'h0888fa08f3f50051fdfefb5ef4af0711fa12;
mem[761] = 144'hf2befe1afa910c440cc70a3208d8fa4f04f5;
mem[762] = 144'hfc9bfa13fb88036cfcfc0f300b20017e0fc2;
mem[763] = 144'h072bfe7f077ff1d8f8f1017500f7f6ce0619;
mem[764] = 144'hf1b90d04f8e5f48bff74f775f1b1f37002be;
mem[765] = 144'h0daff0850a6d0ba300b4f6ee0572076bf4a0;
mem[766] = 144'h012400a00a84087a0b090b2205c20b3cf8e6;
mem[767] = 144'h09a20e4cf03701c5f6d8f17408dc058c04e7;
mem[768] = 144'h0dcbfdedfc08fd9f008bfb9e0f600c98f060;
mem[769] = 144'h0ad20ce60c37ff9efe4afe88082df5bf02d4;
mem[770] = 144'h0e360952f3e8046b0559fc04f7e30e7a07de;
mem[771] = 144'h0f1108290561047ef90208fd06a6fec90db9;
mem[772] = 144'h07eaf20c00480fbdfb4d0290f1d1f053f632;
mem[773] = 144'hf5770651ff200f7601a1f554f5b606fa02b8;
mem[774] = 144'hfdd100eb070bf93303290edc01c0f6aafea2;
mem[775] = 144'h0257f016080f0b19f51bf2df047303dbf334;
mem[776] = 144'h0034f0a6f66301c704f1f8d3008705800f9b;
mem[777] = 144'hfd03066608c3fa54051ff525faa3fbd5fc2c;
mem[778] = 144'h0a92f67c0cb90de501b705e7fb3c0655fb8e;
mem[779] = 144'hf11ffec502d9f22b0652fce6f1cc08800d94;
mem[780] = 144'hff1dfc4af97503f30783fdcaf39df4db01be;
mem[781] = 144'hf1cf0d430b74f829f2850cde0a88f3a5f302;
mem[782] = 144'h0d930b35f9740a61ffb108660cacf3d308f0;
mem[783] = 144'hf0280eaf0529ffedfff3fb040b8c0f9c0198;
mem[784] = 144'hffcb027af715fe83f3f003140ab908b0f2be;
mem[785] = 144'hf676fa68070004ce026600170f9df2b409b1;
mem[786] = 144'h0ce705020859f2e6f97c0964005b0afaf666;
mem[787] = 144'h08bf00d5fe0c0317f03702130849f3c1fd96;
mem[788] = 144'h01620b5908f3ff410848f7ebf6910d990d36;
mem[789] = 144'hfb11f370f9ae09f2f0770bfaf5baf9310c5a;
mem[790] = 144'h02740c58f1720716055ef72ef15af2baf2d8;
mem[791] = 144'h045bf643f5f00fed01eaffa4f6330d09f587;
mem[792] = 144'h0db30a8ff1fd0b300ff10e780096098dfde3;
mem[793] = 144'hfeda037cfaf6f7290a9808f6f851f67df9ba;
mem[794] = 144'hf0aff862f41401d8f8a9fe390d9cf418fa86;
mem[795] = 144'hfd06ff7b05e6f3aef47400e6095bfaf7f4ba;
mem[796] = 144'hf9020e52fc39010b0deffe2df5f601650ebd;
mem[797] = 144'h05620ceef6acf8fd026f0d09f94ffd640350;
mem[798] = 144'h085b0dadf7700b04f85103b6fbebf457f77b;
mem[799] = 144'hf8cbfee10ef2f2fe008a07d0fc12fef5039a;
mem[800] = 144'hf88f04aefca20c6bfbbafde0093202cd06ec;
mem[801] = 144'hfc94f5730e75fbabf0ed07110648f3ef0c26;
mem[802] = 144'h034f0163028af26403270a0107af0deaf127;
mem[803] = 144'h030b0b10f561f528ffdef0bef6c3f505f71b;
mem[804] = 144'h00d30f2ef14b0f71002d0df2fee50d1e05e0;
mem[805] = 144'hfb73f65f030efef70b69074bf49f03120ca7;
mem[806] = 144'hf41909de09900028f2650c16f5190b7af437;
mem[807] = 144'hf6ccfec001f5047df5f8f4b6072f06bd0d5f;
mem[808] = 144'h01750f820c470acbf199f9dc01620983fcb7;
mem[809] = 144'hf6e2fc5af1ca07200b600ed0048cff80f943;
mem[810] = 144'h0f0e0a13026afb01095a09f1054cfb7903c6;
mem[811] = 144'h03670e650b58f1200dbc0eb7ffaff511070d;
mem[812] = 144'h0b0c0e6d0b67f22c0e5408a0036f0b070d43;
mem[813] = 144'hfe84fa3d0b6105b10f2efefe0c1505a0f7e1;
mem[814] = 144'h08def247f170f3660701eff90658fa36f41a;
mem[815] = 144'h0cb3fff2fe6dfcf009d30b81f5bd04bc0271;
mem[816] = 144'h0616fc9d0cc1f068f8a30619ff00f7530f72;
mem[817] = 144'h05ccf6b00f4b0954f016010df1d903eb09be;
mem[818] = 144'h0da3fc5f03e0f5d6f4db0cebf8220f26f609;
mem[819] = 144'hfe5e0a1c0638fd5f0fa1f03d0eeafd6ef45d;
mem[820] = 144'hfd030dba0cd5024e08810210fec0fc3a0c6d;
mem[821] = 144'hfaee0ddff6cbfc2c0300f23cfde8fefa0122;
mem[822] = 144'h029bfa63fc9f05acfc900e4c02c6f0c90248;
mem[823] = 144'hfe4a01d2f1f4f501f3260c04f869f3c2093a;
mem[824] = 144'hf72c0f560761f41cf930f842fefdfb32fca1;
mem[825] = 144'hf239f4410756fb41fb50fc090eebf4d40c5d;
mem[826] = 144'hf3650c120712fdf5f1050d220215f91b0049;
mem[827] = 144'hfe470fd8f19ef9270731ff97fbbdfe70feb9;
mem[828] = 144'h05090f950688f0eb03ad0f8c0f8bfee70846;
mem[829] = 144'h0ecf0beaf0fcf5420e4ffd1703ddfe6207c9;
mem[830] = 144'h08bcfbfef35206fb0a43f0fb08450c3d08a9;
mem[831] = 144'h0cac0ac9f7ef05590b9f0fd503b40a080a87;
mem[832] = 144'hfd460bc90d8efdbd09f70144f07b04430293;
mem[833] = 144'h0da8064df6090ccdff0bf4ee036103070fc2;
mem[834] = 144'hf3be0a4fffadf103fdf6014a0b0ffbeb027b;
mem[835] = 144'hf4e9f4380d97fbcf079d0fa5ff800550f853;
mem[836] = 144'h01d2fd1a076cf770fb990c25fb3b067106cf;
mem[837] = 144'h0d43f66b0632061d0b7af4ba0c27022d0829;
mem[838] = 144'h0571f852f51909a0f742f5f60047f7f703eb;
mem[839] = 144'h06a6f81505d6f0dcf9870c3ef78f0bd508e9;
mem[840] = 144'h05f10336f3d1f80cf502f17b047ff0a2f530;
mem[841] = 144'h071804b0031dfbf6fc9f09b402b00b03f4cf;
mem[842] = 144'h06e7047706ff07a205c7f683f5770c5d022e;
mem[843] = 144'h043ff85ff180f76007ebf35d03e0f8b4f89a;
mem[844] = 144'h0ee6ffea07d7f6130df007150b890022f7a2;
mem[845] = 144'hf29f0293f174fa9df3280f5bff4afb59fac4;
mem[846] = 144'hfa98f589080f09430f98f804f7b00057f00d;
mem[847] = 144'hf306f5f6f463f793f2c7f8610a2302d200aa;
mem[848] = 144'h0d05072e02710dca024b02edf69bf294f1a1;
mem[849] = 144'hfbea0258f5c305f1f363f3e60f9a0c72025b;
mem[850] = 144'hfae7030af70d0732f0670a2b0138fa44041a;
mem[851] = 144'hf6ba083efbcdf291f9f1f673f1ff0f1a0162;
mem[852] = 144'h07610cd903b4f3be0d990fc4fe1c0583ff84;
mem[853] = 144'hf550f11ff948f35408cd0e02ffda0d1dfd37;
mem[854] = 144'h0a92f8a80c8605d40e2703bc0fd0037c0623;
mem[855] = 144'hf05d0fa705590e2bf73504ea0083f1e60be1;
mem[856] = 144'hf8cc025cf617fab30d5af951fc170198fd38;
mem[857] = 144'hf6a201a7f12ef934f1cff49f0b8d00bf0cce;
mem[858] = 144'h0e960d1d06c0f7800bec02aeffadf52a0d03;
mem[859] = 144'hf7f108c30cb90d4cfd12fdc9fde4002808e4;
mem[860] = 144'h0705f0f1f7a2f6b8ff980ae3f9b90fd90687;
mem[861] = 144'h09890515012df77dfd7106e503e702a60842;
mem[862] = 144'hf1faf38f06fdfe3f03000b49003702b10c57;
mem[863] = 144'hf2b7f83801c9f68407050790fd99f1b7052c;
mem[864] = 144'hf7ebf04ff207fc83fd7d0958f981f80904d8;
mem[865] = 144'h0c20f1abfb8403790ed90112f9faff04fff3;
mem[866] = 144'hf12c0903f49cf49cf75406ab0d1f0910fbac;
mem[867] = 144'h066903c00470f78f03360a58f5b5f8f2f2a1;
mem[868] = 144'hf964ff81082af42c0cd50e47fa8af4150aa9;
mem[869] = 144'hf630015bf623f0e8f35b0c30022dfd54f0c5;
mem[870] = 144'h045008560c8ef3b2fb800b9a0f5efefdfd4d;
mem[871] = 144'h01d6fe4af44bf3550363f0dd09e7f00b0d1c;
mem[872] = 144'h0ba0fb81fcb00763f38df3a6f694f7990048;
mem[873] = 144'hf981f978095efac302730c3000b3031b0080;
mem[874] = 144'h0ac002120940f5ad0fbc0ea30e3ffd260526;
mem[875] = 144'hf4be0dc1f24cfbfdf8b50da4066f0cea01a4;
mem[876] = 144'hfa370b53f40afde501c3f3d6f5fdf60df550;
mem[877] = 144'hf6f905e7ffa908d20543f7a9ffe2fe680a9a;
mem[878] = 144'h0d490346fdc9f3900856fdd1f8250f1ff2eb;
mem[879] = 144'hf3770307fa43056a0c28f6b40051f1d1073a;
mem[880] = 144'hfa66fed2f74f069008f806f205630456fa99;
mem[881] = 144'hf503f74402e307900dddffe3f7b704eaf116;
mem[882] = 144'h013a0f9b04530459f870f161fb38f6ca045e;
mem[883] = 144'h0e76fcb60c530fd10903fb81faca01000310;
mem[884] = 144'h091bff07f91a07bd01a7ff4e024ef66ef2e7;
mem[885] = 144'h0eb5eff0fa1ff639fc68fa2ef29bf2a1f635;
mem[886] = 144'hf68e0f1d0ad10e87f91bf9ac0846076ef436;
mem[887] = 144'h0152f18b0c5f01c5ff150e71fd59f99b0d8c;
mem[888] = 144'hf8ad0bb0070405acf21c07a2f107fb6df8ce;
mem[889] = 144'h0239f161094c0a84074bffa9fd00f9d2fa97;
mem[890] = 144'hfc9d0239ffb8f508097df8ca05c706710928;
mem[891] = 144'heff4f63ffbc503cef8c40e0af19efe0d059c;
mem[892] = 144'h0f13f00ff99f0024f97cf6030d1df8bcfb6a;
mem[893] = 144'hf7e105c7fb47fdb109aef64108b7064d07d8;
mem[894] = 144'hf1610717f3a10919f4b6087cf08400fff018;
mem[895] = 144'h0ef3fef20bac0a2d0b8a017b07100f28f2f9;
mem[896] = 144'hf9a803830300fb560999f26808a0f882f645;
mem[897] = 144'h01c90b9b0d93086c00d4f95ef5ff00ae0993;
mem[898] = 144'h0791092d09ab0946005df4aa0dec0eaf0c83;
mem[899] = 144'h04240ac2ff670d19f390febd0c240dbcf0e2;
mem[900] = 144'hf26df55ef699f46d00acf3ff0fc10ce3f0d0;
mem[901] = 144'hfe8402380dbcf84d0f02fe97fdfb085cf71b;
mem[902] = 144'h0cc1045302f2faa0f2d7f541f742f608f9bb;
mem[903] = 144'hf0210627f54f08450d80047003d7fc75fcb7;
mem[904] = 144'h044f0a32fbe2fa540468f8330c89fd4c04ae;
mem[905] = 144'h0822066f0d430d930cedf4c4010efabff162;
mem[906] = 144'h08ee0768fbb7074804c7fb520bc0fc7df8a8;
mem[907] = 144'hf0130f9af37bff860a75f249f5fa0a490756;
mem[908] = 144'h016608260aa9f0920adb07b2f84dfbf9f2b5;
mem[909] = 144'hf3bfff6df9fffc0b0b5505ec0ea8efdffa3b;
mem[910] = 144'hf7ec010cfc980e7505d5fb7f0ba1fec60928;
mem[911] = 144'hfff40a7606cef31200bdf38cf47d09a8f0cc;
mem[912] = 144'h0c13f3d5070f0f93077b021dfd2c0eb9f36b;
mem[913] = 144'h0e6efb5ef00a08d5f7110acafea6087a0c42;
mem[914] = 144'hf5a40b480562021df6d7f7540da40dabf812;
mem[915] = 144'h0c47f13103f0094e0286f34bf12cf522fe82;
mem[916] = 144'hff18f2a604def5fbf5b8f20c06f80c89fabe;
mem[917] = 144'h0741fe1305220f5d001606ae0646fbc601ca;
mem[918] = 144'hfc810ae0fd21f9f9045a06a30726015106b5;
mem[919] = 144'hfe68f773012d0109fd92f298f57bf8e7f904;
mem[920] = 144'h0058f8a0f8e4fb4ffe930a77f145041003c1;
mem[921] = 144'h0a02f3cb01c104e4ffa8057cf8ecfe780aa2;
mem[922] = 144'hfedbf39b0921059d00f50de00f160a88f5ce;
mem[923] = 144'hfa7208f305ed068df65309170c7af093fa8b;
mem[924] = 144'h00fcf857fed706240034fcb60539f12ef6ae;
mem[925] = 144'hfc74f823fc6f045b0827f27309cf00e209bd;
mem[926] = 144'hf94f074aff8a08990a69064b04f0fdabfea6;
mem[927] = 144'h0d3ff18af04beff00bf40fa8ffee0398ffcf;
mem[928] = 144'hfc9ef0910d42f3bbfa250002f6b606d2011a;
mem[929] = 144'hf10d05ff0d5e0bbe07b3f352f6d2f29c01b2;
mem[930] = 144'hfda1ff80ff15fc13fafbf7be02cafbb1f926;
mem[931] = 144'hf6e9f301fed0f4530bd808f9fb5c0916fa87;
mem[932] = 144'hfcc504420db3fcaf037cfc5ffb8dfc15ff94;
mem[933] = 144'hf2be0b0807e4f663fc64fd8f0f4fff7df241;
mem[934] = 144'h0c620b1901c30528ffa602a40544fe77f69c;
mem[935] = 144'hfaa2f98cf116fefc0368f8f804fc04a80886;
mem[936] = 144'h06c3ff1ff357fa53fc9e0831f9430aec068a;
mem[937] = 144'hff820caaf44d0976fac9039305aef1fb0d5b;
mem[938] = 144'hfa45fb2df2ccf186f92701d3fdd10b710ac6;
mem[939] = 144'hfd2e00dd0d6c0e4afc3404d701bdf16cf419;
mem[940] = 144'h0a3a0c37f682f49cfc94fd7df8ddf398f7a2;
mem[941] = 144'h099ef632f77006a30abb0c3dfdd00110fda2;
mem[942] = 144'hf1a60f33ffb8f3190857f7620c55f6d1ffed;
mem[943] = 144'hfb62fc4b042ff2e2f95909adf738f880fcab;
mem[944] = 144'hf48bf27ffec0fa00fca7ffddf1cffb3cf027;
mem[945] = 144'hfd0500c3f592fd310c03f51bf9b2f7a5f66b;
mem[946] = 144'hf31e0bec0e320a4a07ecf570f33dfb01f3fc;
mem[947] = 144'h05c40e1bf349019c0612fe75045ff3150e1c;
mem[948] = 144'h0d27f9f309bffabf074701d30253f801f736;
mem[949] = 144'hf6b602bf0ee6f17b018800eafb39f923fd3b;
mem[950] = 144'h021001870129f484f84afe59039e0ed20740;
mem[951] = 144'hfae2f7f509d40668f233084ef943f8170df8;
mem[952] = 144'hff64f1df0943fec309b2f7ebf1bd0ba6f7e7;
mem[953] = 144'hfecef18bfa85f90af7eb032ffcc9f9320dde;
mem[954] = 144'hf764ff81fd630650f3120420091c0649f18d;
mem[955] = 144'h0b360513f8c7f5e10dda0ce7f76104adf275;
mem[956] = 144'hfd7cfe6301b60f8004f9ff6ff41dff84f7a8;
mem[957] = 144'hf078ff40047c0d3407f3fbbcf8ec078a0038;
mem[958] = 144'h0a44f894fa1af1ecf0c9f8be0dd1059ff0b0;
mem[959] = 144'hf07df328fc92f83007f6ff8af601effdff59;
mem[960] = 144'hf5520277f54a08affbeb0bacfa75f8e4f22d;
mem[961] = 144'h00a3f985f0d4fc44f6e60061fce3fed2010d;
mem[962] = 144'hf9affaac02ecf9c1fd3cf785fbbd062900e6;
mem[963] = 144'hfa08fca8f38ff1b9f7c6f9810a7d0c40f9aa;
mem[964] = 144'hfdb2feecfb36fead0c070d84fc2b034901c0;
mem[965] = 144'h022cf193fd92f2bf0f2b0e52f39703810270;
mem[966] = 144'hf05bf7eb06d1f8e10761fe610b34fa35fc5b;
mem[967] = 144'hfde5f2b802f4f8c4f0b8f6200f7c0f61f8d2;
mem[968] = 144'hf714f03b00420bd7f1e30608f2e20e36ff98;
mem[969] = 144'hffdff84b023e0f4f0b6a0891f43605f8f9a0;
mem[970] = 144'hf556f39d0ff9f09c02dd0a53031cfa08f42d;
mem[971] = 144'h03b4f3e3024102cf0f760c2201b10b190923;
mem[972] = 144'h0fcefb3508130eb0f1ae0b68f298f9c30392;
mem[973] = 144'h099f0f95f4d6f9dd021404ce095b0c5df489;
mem[974] = 144'hfdd90644f543f808f7390826fdc10d7c0912;
mem[975] = 144'h0abb0e44f86afbcf0d280284fd9df347feea;
mem[976] = 144'hf2b309f2fb070d34fd47f0b40bb0f054f8dc;
mem[977] = 144'hf4f2fe2cfea70bcefd59f4ddfc0bff1e0116;
mem[978] = 144'h08f6f691f741fa38f1c8f8d0f8d306ee0a43;
mem[979] = 144'hf0c80108f37305a6faf7fb5ff16d00b6fdb4;
mem[980] = 144'h0e3ef6c1f8a5f34bff250de5fbe8040305cb;
mem[981] = 144'hfa550600f9affb6ffe50ffedf8520b2c0ae9;
mem[982] = 144'h0143fc0dfbed05190e52f3c4018bf67bf0ac;
mem[983] = 144'hfc310226fcfbff02f442f0cafe680587fbde;
mem[984] = 144'hfd1e0ae003500e6ff21df30e0eaa0c89fa4c;
mem[985] = 144'h0840f27ef6eb0ddf01cef8bd029df4abfb9a;
mem[986] = 144'hf47e0786029409f50d420ca204f10b30f989;
mem[987] = 144'h0707f4b3fc9407cbfbdaf55e0ec1fa8c0094;
mem[988] = 144'hf4f2063a06fffd37fffb0674fdeaf70bf311;
mem[989] = 144'hfc91fe7efaebfbee032ffe95f152f80b0d9b;
mem[990] = 144'hf0a302960e6ceffefc79f33b00f1f8b3fe55;
mem[991] = 144'h0b0a0868f74d0cccf7cc0ebefcdff386fd84;
mem[992] = 144'hf2830beb09f7f022f0b30f89039909350f7f;
mem[993] = 144'hf51b034b0dcdf146ffeff76e0c82f9d1f4fa;
mem[994] = 144'h0124ffbe05df091efc7b0e71f87f0997f995;
mem[995] = 144'h0a070cb4fe400a500173ff5f09160f060522;
mem[996] = 144'hfcf1f00b07d3f573080d0a5ffd93f0a10ab7;
mem[997] = 144'h0e60f3e50b540a9a0b900a010fa20441058c;
mem[998] = 144'h0ab8012df7ac01340ec5efd00ca101fd04cb;
mem[999] = 144'h03d8f84a046b0b6ff488f3fcfb010527f889;
mem[1000] = 144'hf897f2e8f18201e70e5306b800b4f39904a4;
mem[1001] = 144'hf9210d9a07e6f7e10eca0efdf3b90f18f99e;
mem[1002] = 144'h0105015c085c0277fbd6fcb0f1e10bdf021d;
mem[1003] = 144'h071a09c8fe58fa0bf02f0741f77a092808f2;
mem[1004] = 144'h02da0b7a074ef7d409f9f161fa04f0f5f2c5;
mem[1005] = 144'h0e8f0d8c0b430ca3f3d9fba9f5620877feb3;
mem[1006] = 144'hf7aa0f2e00dc031a0958fc70f9ddf07906bb;
mem[1007] = 144'h04de00c8ff29f0b3f70807e407bc03440bba;
mem[1008] = 144'hf51b0ae6f48eff080783f726073b0f53fc69;
mem[1009] = 144'h0dd0fec4f5530c7b04a30cc90ec2f003faf4;
mem[1010] = 144'h089cf0fffa42001eff2efb16f73f02ff0934;
mem[1011] = 144'hfdb1fada0de40d2af229fdccf19e081cfc2e;
mem[1012] = 144'hf7c2098607220486f5cbf5df07c70a3b0caa;
mem[1013] = 144'h02b80de7fc7bf0c0f45907520a93ffba09e2;
mem[1014] = 144'hf6e6f136052bf8ee0a490cb6f057ff3c0424;
mem[1015] = 144'h069df0dcfb81029bff02faf2027e0909feee;
mem[1016] = 144'hfaa9fff4fd3c0e0e023e045f0b2606b80f4a;
mem[1017] = 144'h09d4f00305a1063d0d7cfe480deb0f76fc7f;
mem[1018] = 144'hf005f420fbf20c42f912fea2fb66f7fffe37;
mem[1019] = 144'h087a012e0c39072bf3f7f5f0f03df8010d42;
mem[1020] = 144'h020a052b07e3ff5f0b66ff25f7aaf057f645;
mem[1021] = 144'h0e11fe7e0d1d06a6fa7a0118fc2cf3f1f86c;
mem[1022] = 144'h0121fa27076e048af5fef89a06010386f2c1;
mem[1023] = 144'h028d07cafb090fcc027bfa040274f597078b;
mem[1024] = 144'h0d3d023e080409a3026d0cc6f879f26702e4;
mem[1025] = 144'h04c7feb2faf00f610d67fb08f95c09a6f14d;
mem[1026] = 144'h04720a7b07f7f85a0a66f97ef00af31cfdfc;
mem[1027] = 144'hf2d70521043af4b5fd22065cf97c0700f43d;
mem[1028] = 144'h0becfbc70b6a0934f0aefc94fb850093fe00;
mem[1029] = 144'hf3dcf128074ff41ff2f0f4fa07ec0d49f238;
mem[1030] = 144'h0481faa9f0f70f1df5f2f51b02bbf92a06c6;
mem[1031] = 144'hf7a804780ffe0f91fd1d06110c48f2250eae;
mem[1032] = 144'h062f0aa50ab60a880f950c3e03b7046908cf;
mem[1033] = 144'h0684f4070088f73dfd1efdb4fa42f492f4ee;
mem[1034] = 144'hf214f1ae01a5f4fef71eff4ffec20e130da1;
mem[1035] = 144'hf96a0b7e0be3042303a400b2fdd4fb5809ca;
mem[1036] = 144'hf91c0404fe5d0e1d094e0afc0d7cfa6b07cb;
mem[1037] = 144'h0f41fa2b0f900e230ef3034d0a58f1060952;
mem[1038] = 144'h0d510e6f003801ab007405590e8df0f10ece;
mem[1039] = 144'h0870fea0f912fba80099f3620dda015e0c67;
mem[1040] = 144'hf7570dc008c2073f0c6dfef5f418fef302c5;
mem[1041] = 144'hf3b00285fee2f24afaec015df482f94e0478;
mem[1042] = 144'h0c8ff86e0fed076ff9b6fcef0c9001e3019b;
mem[1043] = 144'h0db507420dbaf9c1f7980563f8a7f012f312;
mem[1044] = 144'hffcef07c0d66fbe9f4200d34040c0d1afcc9;
mem[1045] = 144'hf89a068c047af5cdfaf5093f086ffb180235;
mem[1046] = 144'h06a70992fc52023908e30ae3f8f0fcee0984;
mem[1047] = 144'h061c031d068b0df208bff2e009def7b6f328;
mem[1048] = 144'h06fc04d3fc95f885f5f1fba10872f22cfc7c;
mem[1049] = 144'heff80feb0469065ef251ffef070cfd7bf51c;
mem[1050] = 144'h0b3ff3550cff0167f1a7fcc2facff0970ff7;
mem[1051] = 144'h0f92f47b0d910cb6f95cfe97f0fc0e5ff3a2;
mem[1052] = 144'h0c56fef0f71bf61908480e13f5bfffdf0782;
mem[1053] = 144'hf6190a58fa9bfb340043f4fb078ffcccf1d9;
mem[1054] = 144'hf0a6f1660be9f787fbc8ffbf05ba0c68f7a6;
mem[1055] = 144'h08f7f03ffcde086b0048f64af9c6022801bf;
mem[1056] = 144'h084aff5bfe080844fa76021a0eedf12efaac;
mem[1057] = 144'h04d1fd820a8cfa65f2d802d80fa605390f2a;
mem[1058] = 144'hf1f0059ef8a1f5360a4cf9aafe83f1600f8e;
mem[1059] = 144'hfc81f6ecf1e108f4ffa5f0380d3bf66bf9a0;
mem[1060] = 144'hfd8d06e1f89bf9cf0b8501170b4af3cbfe15;
mem[1061] = 144'hf4a708490b780e3af23ff05f0f17f079f32b;
mem[1062] = 144'hfa98ff8f08d60711fe8cff3e07a7ffdb058e;
mem[1063] = 144'hf629f610f6470e3402c1ffe405b5001d012a;
mem[1064] = 144'h02c6039dfcf1faa00e5bf530f2c2089afe69;
mem[1065] = 144'hf4fcfa240e29fbd90f12f1d10a6f05fa0b42;
mem[1066] = 144'h031ff1ff0d10fc5d0cbc0af8f131f461033d;
mem[1067] = 144'h0ed8f246fb40fd3609f50eda0162ff660ecb;
mem[1068] = 144'h009df2c50dabf216f6b80c73001608d9fe73;
mem[1069] = 144'h06d402c2f1bc02fefa3b09f403f2f552f4d4;
mem[1070] = 144'h0b12f1c302d2f627fcc9f4ca09e3f932017d;
mem[1071] = 144'h0f1a02220d95fcebfbc2002605d8f773022f;
mem[1072] = 144'hffde0bd2f2f7fca3044d0acffc6e00120480;
mem[1073] = 144'hfea8f788f53001b4fc78f9e60933f4610007;
mem[1074] = 144'hf59f09670dd10d79021a083b0282083e0612;
mem[1075] = 144'h02d001c6f9d2ff9709cbf287035ff8540a5d;
mem[1076] = 144'h01acf6fe06050cb9097efe72f3d70e46f9e8;
mem[1077] = 144'h06f30669fc7e0fe6016c07250c44f18b06e5;
mem[1078] = 144'hf180f834faf50c23f403fa15f6db093ff8db;
mem[1079] = 144'hfded05f20a84021df6f9f4280fbd0ba8f9cd;
mem[1080] = 144'hf2020595f8fcf55b04a8f5b9fd04fa0501a8;
mem[1081] = 144'h0502f0a4f0ca086ffbe3fe1ef1f7033b0899;
mem[1082] = 144'hfcaafb87fe7bfc76f661fae7fcd3f54609f4;
mem[1083] = 144'h0d51f5c70b6af929f639029e0352f569f088;
mem[1084] = 144'hfb2d05f00fc3f67f0ab70e35032bfaa10b34;
mem[1085] = 144'hf86af3a3f18eff4401b1f8b0f4800a0d0460;
mem[1086] = 144'h0d52f3ab02a109a1fa02f7280c86f18af416;
mem[1087] = 144'hfc1afcf6f51a0c38034bf0d9ff68f817fb55;
mem[1088] = 144'h0cc00683fc6c09750151006bf7730656f4f9;
mem[1089] = 144'h09050c880e66f6a2f6aaf5dcf59df21108cd;
mem[1090] = 144'hfb96ffcc0364fcb008a00a8a0cd3f270fa9c;
mem[1091] = 144'hf188fcb3f056f99c0cbf01981032f72e0451;
mem[1092] = 144'h010cf66efb6d0d8cffb00ea9f21afb790f9e;
mem[1093] = 144'h0943f20afe050a90f57d08a60fa6fa640038;
mem[1094] = 144'hf0b7f9df0de50049fafdf634fadc058bf5aa;
mem[1095] = 144'hf690fc92f927fa40f9550422f505f308f829;
mem[1096] = 144'h0ad90827f61ff88a07bd04bcf34e06140b3b;
mem[1097] = 144'h0bfbf5bf07c6f91f0364f8def6be031b0bff;
mem[1098] = 144'hf4aaf350f38d0f5ef91205c80301fc7af94e;
mem[1099] = 144'hf6c70a05f94804fa01aefadc0e3f0023fe85;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule