`timescale 1ns/1ns

module wt_fc1_mem4 #(parameter ADDR_WIDTH = 10, DATA_WIDTH = 144, DEPTH = 1024) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h0f000b9b0062f92d0ac6033f0903f404f12e;
mem[1] = 144'h040f0491ff8006f40433f99afbedf1fff1f1;
mem[2] = 144'hfe49ffcc09040f300c1b03890007f1cd0d86;
mem[3] = 144'hf9faf0a00702f92ffea7f9d0fb58ff19f04b;
mem[4] = 144'h04b3f9f4f84c0920f66308c3fdf802cc015b;
mem[5] = 144'hf4b20c15f171094d0c6108eb09440aeefdb0;
mem[6] = 144'h05620327f2ce0ddafb1ff58cf14ef1bef704;
mem[7] = 144'hffb9f54df3790ddc07ae0101f33df9aa08ff;
mem[8] = 144'h0a02f8c7037ff29cf7420e42f09cf93807af;
mem[9] = 144'hf2d7f82f041107df029400f006ac0e7d0acb;
mem[10] = 144'hf5b1f6f0f0c8f7b7f3020ee9f6fc0021fdd3;
mem[11] = 144'h017cf2fc001b0aef01490dbb026608bf0734;
mem[12] = 144'hf02ef9b2f067f1d4f6b90c11f3ca07bdff47;
mem[13] = 144'h0aa70b04fef90a96f369fd3608d0f01002a8;
mem[14] = 144'h051cff0305ba02a0005001cd0306f33a096c;
mem[15] = 144'hf3c401bdf920fc71f579f0f0f69df6ba0604;
mem[16] = 144'hf312fdebfc650d940885036ffddff150f8ea;
mem[17] = 144'hf6970927007d088ff4b102a7f84d05b005fd;
mem[18] = 144'h0edc00fef54b0d81003affafff510887f858;
mem[19] = 144'h0605f7450525f8a4022a0270f47c06fb0a96;
mem[20] = 144'h0875f2d0f017f9b304f0f015f6f203cef78a;
mem[21] = 144'hfd850606f95efc61f19c0f0c0013f0e4fbaa;
mem[22] = 144'h0927f1fcf6def99109e50025ff3505f8f6c9;
mem[23] = 144'h0ff9f4b7ff33f50ff4a30bb80293f7abf962;
mem[24] = 144'hf1f8061ff465f022f856f4bdfb9ff76801fe;
mem[25] = 144'h0cedf16b026dfb9a0bd5fe240ae2f0d00cf0;
mem[26] = 144'h0e4009b2f60a02f7feb3f66e043ff55805a5;
mem[27] = 144'h0bf7fceb0d8af11f051afaf4067ff517f473;
mem[28] = 144'h0e240c0bf6000f88f9810f44fd55fcfdf1ec;
mem[29] = 144'h0777f9b0f5c9f0ca02730510f527f74ff7be;
mem[30] = 144'h0700097902040ab400640a140d810ce5f012;
mem[31] = 144'hfe4600d2f7fc046c00cefc12f5650378f064;
mem[32] = 144'h0bf7eb24ff0bebeeede5fefbf449eb1ce1a6;
mem[33] = 144'h0f5bffab0ab20d7e01bcf35b0a5300b10487;
mem[34] = 144'hfe92f0d1ffbbfe68f075fde4024f0640f713;
mem[35] = 144'h0ac3f9c4fda8fb15f47ce406f154ec12e56a;
mem[36] = 144'hf7f1f514f736ec76f5f00132069c00c7f103;
mem[37] = 144'hf978071b0dfa01a9fe2df9e0f5b70593f39e;
mem[38] = 144'hfcfdf823f27d0ca5064300ff064106da08e6;
mem[39] = 144'hfd0906cd0b01f3b5004bf9c1f14ff3bef510;
mem[40] = 144'hf626f050049a0c73ffd3fb53f0cf01400263;
mem[41] = 144'h0479fe7701e3f219f50b033e0050efadfa2b;
mem[42] = 144'heae6f68d07670650f645e486ebdcfd35ff96;
mem[43] = 144'hf65505e2f3d7f9bbf3b3ef02f6f70a8f097e;
mem[44] = 144'h009304d4f4f9f37001bee73703d2ef7ee378;
mem[45] = 144'hf5c7f673f31ef005086df76d0f5ef1d4f477;
mem[46] = 144'hf830f018fbc6f76cfafa0b43f125e293faa0;
mem[47] = 144'h006a08e807c209ab09d6058a0c1503b0feb7;
mem[48] = 144'hf15beabef076fd72f2250310ea3ff448f6ad;
mem[49] = 144'hfde7fcbbfd2207f1fc910971f1e1ff570882;
mem[50] = 144'hffc007c3f83df67308d4fc910ee406bf06a2;
mem[51] = 144'heef3f702f83cfa18eed0011eeb34f4fff7e2;
mem[52] = 144'h08920829016f05d909c9faa407b3f075f760;
mem[53] = 144'h00d3ff2ef5fbf98508b90b750826f49a073f;
mem[54] = 144'h061306100882fb760f2701220636f3590d71;
mem[55] = 144'h077c0b5006f0fb9809e1f02c0bfafac0f433;
mem[56] = 144'hfadff8cffcc4061c0d74fc9ef37cf999f2b0;
mem[57] = 144'hfa21f9660426fb57ff420f13f48605b60255;
mem[58] = 144'hef95f7c8f416ea09f6a4fa5be05ee6fa03e5;
mem[59] = 144'hf3ff04db09ee040ffcabf0f70cb907faf0c8;
mem[60] = 144'hf56505b602b9e8c4f391f28aff00f910ecf5;
mem[61] = 144'hf457f2b206e9fb1407de0afef5d7f8d00155;
mem[62] = 144'hfe280484fe4b02aafa12f069f730f7d5e880;
mem[63] = 144'hfe6af956f1cbf61bfb8601140680ebf3f61c;
mem[64] = 144'hf2c3f941fb5df1da03b006ff01fd009c0552;
mem[65] = 144'h0a8d0b95fc74fa81f18d0bebf82af6f10147;
mem[66] = 144'hf06e07f4033afb81fb0af470fa01f4c2fb8f;
mem[67] = 144'hfbb6fd2aff94019af77ded7ff8d5fa9ff88a;
mem[68] = 144'hefa100b9fca5f621facefa810275f27eefad;
mem[69] = 144'hf418ef95f0cafd4ffcaaf3b0f0e7053bfea4;
mem[70] = 144'hf8da0dc4028100ee0d88fd3c02190c79f6e4;
mem[71] = 144'h0ca2fea002030807f681f55ff78701d3f31a;
mem[72] = 144'hf650ee9a03d205a20bdd01ef0ac800ccfd70;
mem[73] = 144'h04d2fc4aff510658ffd9f628f117fc79f15f;
mem[74] = 144'hfceeec96e89df1b8eb74f461e2e8fd7f078a;
mem[75] = 144'h0678ef3e0aa3f123f5b2f312f6dcf976fe9c;
mem[76] = 144'hfe7afae6005de580e5e9ecaefdc2ff18f199;
mem[77] = 144'h04f902ba070bf682fae1f60f02cd09cbf196;
mem[78] = 144'h09b5071502590527049b0714057bf9c6e0d0;
mem[79] = 144'hf7f20bbcfcd9ff27fd93f7c6fb6300eb00d2;
mem[80] = 144'h032df7aefbaef498fc0afd0ef0b2f10ff153;
mem[81] = 144'h014006a60e770c2af45404b801ab0af60a8e;
mem[82] = 144'hf625029ffe9407c70b260bd8f818f9b30b4b;
mem[83] = 144'hf9b905b90206f7aef64df2110caef235e955;
mem[84] = 144'h0b92fd4d094d0c500660fc7af2cb01fff30d;
mem[85] = 144'hf62b013ffa3afb9a00a209f00ecc03be0ba0;
mem[86] = 144'hf45bfa4bfa160374f2e601c8fc4bf25a0ab8;
mem[87] = 144'hffe0ff820fc40e55f57e0d1efece07dc0842;
mem[88] = 144'hf6bbf1f9fa70f383f3e7fd69f982f2b8feda;
mem[89] = 144'h0444f992f2a40af00a7e06840bfd076c0767;
mem[90] = 144'h0763fe39f2140db3ffd7ef79fa2f0764fed6;
mem[91] = 144'hf8fbf17d02e80b4c03cc04b2ff44095def70;
mem[92] = 144'hfbf4fd7dfc6ef3c8f50df705fe0ceefe026e;
mem[93] = 144'h076efab4f3520ad1fdb8097f015d08d7f420;
mem[94] = 144'h0059efd302a708020cb404560aaaffc9f899;
mem[95] = 144'h01fdeed1f5eaf83af4e4072cf37af2b8f8ea;
mem[96] = 144'hfb4bfad203810146f33a031fee10fe6ff2d3;
mem[97] = 144'hf0c60a5dfab100c7fc6bf1b3036a0a3bf15f;
mem[98] = 144'h0cb9fbd7f82c0cd5fddbff8902c102f4fe6f;
mem[99] = 144'h081fff6409330a61f70808470afc06cc090e;
mem[100] = 144'h0ef7fd1ef144ef2af7fafd41f186faac0b9d;
mem[101] = 144'h0166f508f97df3c8fe21f8f806fcf3a20710;
mem[102] = 144'hf057fcfc03d5fd8df43d059cf14ff29bf04d;
mem[103] = 144'h026b00830bb30aaef99f0ca606b7fe7dffcd;
mem[104] = 144'hfa63f667ff3705faf4be0caefa5008670cd5;
mem[105] = 144'hf573f0b400a2f91c0cccfd010418fae10a30;
mem[106] = 144'h0c5c091bfd0df260fd04020d07ff04faf95b;
mem[107] = 144'h05f5020c0b6efe34f25ff553000609c805a5;
mem[108] = 144'h022e0809024c04adfaadf4f3035c09610f10;
mem[109] = 144'h01040524f581f7fff938015cf104fdfdff3a;
mem[110] = 144'h0a78f19ef14cf857fee1fc8cf4850466f3af;
mem[111] = 144'h015001ee0723f35f0260fe98fde1f111f7f1;
mem[112] = 144'hfa09fd4aff22ed7903cefd9df81ffffb0253;
mem[113] = 144'hf016f018f438f864fe6b0ddffca1ef2507ce;
mem[114] = 144'hfc4aff8b00f70b71034f0b6806f50d3dfe56;
mem[115] = 144'h0760fe2af3b6e74406e8ed5a019aea66ed54;
mem[116] = 144'hfb94fd550bc3fc60f9c20943f09bfb2805c6;
mem[117] = 144'h0bb5fd370233f301f1fcf104fea7f38c0769;
mem[118] = 144'hf0f404f60c2ff3caf18d0053024a0873f312;
mem[119] = 144'h0787fb19f141f208f2ef0adb008ceed50531;
mem[120] = 144'hf8580bea045f050cf63cefbbfe46ebe7e935;
mem[121] = 144'h06d4f2bbf7e80476ef5e0768047dfc990acb;
mem[122] = 144'h0cd8f69dfb00f38afdc2ec90ef77f501f95a;
mem[123] = 144'hf5bbf67803f4060b060f0d57f8a4f447f623;
mem[124] = 144'hf2f8fd8506760274fb6cf3a9fbbcfcc2ff9d;
mem[125] = 144'hfe69f390f80506c7fffe0e20f0cefca80e4b;
mem[126] = 144'h05d5fc070b8b06faf662f100f29a0a1af9ad;
mem[127] = 144'h0ca7ff8704100c2f0846020b0ba4ef4e054b;
mem[128] = 144'h096d0075f8e7f46003e3f3e60e1cfa6afee8;
mem[129] = 144'h0920f30c063ff55cfa96f1d8f83bff240597;
mem[130] = 144'hf34100def2ee0f25fc15074cf296fe6ffbef;
mem[131] = 144'h0503030f09cb0572049d02a3fca60ab2f450;
mem[132] = 144'hf86dfa7bf425f459f8ed072ff62cf6380c08;
mem[133] = 144'h06550e5afd23f09cf7fdf606ff2f0f19039b;
mem[134] = 144'hfb40f026f83604d6039d0212f8d8f3a00af8;
mem[135] = 144'h0ad2f64af5a80389fb1df840f66f0c23fd74;
mem[136] = 144'h076d05ef0f84fbd809860598063d02f0f292;
mem[137] = 144'h05d002640e560e99f6cb0566054d03570daa;
mem[138] = 144'h017308b7f05c029ff9210457073af73ef3b6;
mem[139] = 144'h0352f3850efd05bbf38df2a5ff1403eb0ee7;
mem[140] = 144'hfad00f33001d0c25f566f825f08df644fe76;
mem[141] = 144'h038bf7010833f551063303f7089ef7ce01d6;
mem[142] = 144'hf6450063f6ccfe17f101fd7af0f20656f9c8;
mem[143] = 144'h0947f645f9d4fc05fd9f0401fc79f91bf32f;
mem[144] = 144'hf9a0f951f4a4f2d10d03fb2f0534f1b405b1;
mem[145] = 144'hfe4c013b0d6ff1510b5bf7d6fd2d0e050be3;
mem[146] = 144'hfb23fe4d01f4f4d607140154fbeeff8ffc31;
mem[147] = 144'hfc1b01800e0906d5fbc505e2f012fe7f07c2;
mem[148] = 144'hf821f544026af89e01b90cd8fd8308410941;
mem[149] = 144'h0c2af32301e7fe5bfdf4057df82207fa0517;
mem[150] = 144'h09b3fdb3fc4508750a5df2eef9c1efe3f9d9;
mem[151] = 144'h04b2fa2f07d4f628012cf6a6ffb2fb75091c;
mem[152] = 144'h066dfb7409f401aafffc0dcefb0cf902041a;
mem[153] = 144'hf5b5fd01f208027df7f8f57ff22df6cef902;
mem[154] = 144'hf305f487f83af2c1026cff52f4a4fff5ffa8;
mem[155] = 144'h0421f51ffb47f05ef2d3f74ef0370eb20a24;
mem[156] = 144'hf64504a0f6730b8df17efeb8fea6f4f0f766;
mem[157] = 144'h057e0317f44ef822f44b09a4f6fff53affca;
mem[158] = 144'hf1750b800828f4620782fb4ef9d406dd0ba9;
mem[159] = 144'hf282f13bfa69f116f694feb4fb18f6af07f6;
mem[160] = 144'h0370ff470747f9e70362017efc54fdb70502;
mem[161] = 144'hf93d0b66ff99f576036dfc00fc39feabfa92;
mem[162] = 144'hf5b6f48e0b45f3f0fa1e042ff2c60f0cfe9e;
mem[163] = 144'hf794ff2bf732fb78f2cd0c5c08adf2e2f2ed;
mem[164] = 144'hfad8f38cfbcc00e0fbd408f9fa1d0379f246;
mem[165] = 144'h07c00ee0ff1100caf5e6058a0ec70adf0f22;
mem[166] = 144'hfdf00366f64a00c60305ff0b0077f08a019c;
mem[167] = 144'hfe5a091cf03102d4f2d8fb240540fdad0dda;
mem[168] = 144'hf92d0fc00fddfbe00f380455f7ecf513fe88;
mem[169] = 144'hf31af763f626f03a04a7ff76fe120583f3be;
mem[170] = 144'h097ef965f815ef7afc3dfb69f554ff550678;
mem[171] = 144'h00a7040a0952f0080ce9f394fe41fca8f246;
mem[172] = 144'hf79b0450064e030df3810646f5c7fb410a6b;
mem[173] = 144'hfe0ffb60f38bf160043c0f36f8a8008ffbfd;
mem[174] = 144'h0aaff90d0f5afd48f1080f8b0b7ef32cfaf2;
mem[175] = 144'h0872f4a1f3ccf4f50e7cfe51f53cf496fb97;
mem[176] = 144'hfec8f031f12409f2ff84f4110b60f0c0fcfa;
mem[177] = 144'h0b9ff874002d0d9df64bfd39f30d0b26008d;
mem[178] = 144'hf7f804e30747f6330e61f89cfa2c086106f0;
mem[179] = 144'hf3cefab1fcf40442f942f90806120228fed3;
mem[180] = 144'h0923027cfc34fa6cf3eafa6a0476f6eff4e6;
mem[181] = 144'hfe2c0b5906240117048a0299fa19fb81f012;
mem[182] = 144'hf49d0c640a2003b3fb7bf55ffaf2020f099c;
mem[183] = 144'hf95ff1f607f10d930473fdcef3b9f685ff61;
mem[184] = 144'hf024f20a0edf035ff2eb024c0b46f060fa93;
mem[185] = 144'hf5f1fc1b092ef9bf0e7a0b60fb410cf6f7d5;
mem[186] = 144'h088ff85f08be0d89085b0107f51609a5fd50;
mem[187] = 144'hf9c5f872fb3ff98a00640f23f44005330244;
mem[188] = 144'hf8880b9b097efec205e2f7f306ae0d7a0500;
mem[189] = 144'hff06fe3500c60dd905a4f3f7f854f5530bcd;
mem[190] = 144'hf30707c2f4dc0d3af511f97efaa504b20af5;
mem[191] = 144'h04ecf02209d2fb49fdef07d5021f0234069a;
mem[192] = 144'hf93ff54e0981005c0271f29b028e035e04aa;
mem[193] = 144'h04fb08c7f019f36ef48af538f3e70106fe41;
mem[194] = 144'h04790594013df83e0b3002edfe4c0f310741;
mem[195] = 144'hf54607ac0d46ee14ef1e0a5dede4efac02e8;
mem[196] = 144'h0309f9e907aa0884f455f64e04ccf012ee4b;
mem[197] = 144'hf2d3f0a60c8cf080f70af3effc08030af4eb;
mem[198] = 144'hf9ed02b0f1bbfa170f06071008ed0e53f05a;
mem[199] = 144'hf2df033806b4fce80074031ef6d80606fb0c;
mem[200] = 144'hf9a8002a03300602fa4000020af4083dfdc1;
mem[201] = 144'h0c360460f2cafd1409aafeddf8430ed10813;
mem[202] = 144'h06bafbfa000b008bfebbf84e04b200c806e6;
mem[203] = 144'hfabbf53909050d750148f8950e110671f9a8;
mem[204] = 144'hfef8f0a90335eedbfbeaf9b8f826fbc3f204;
mem[205] = 144'h0e770ff109b3f34afba70dd6f551f47505f1;
mem[206] = 144'hff180ebff4c2fd2bf078fa3bfc490952fd57;
mem[207] = 144'h0c3d021efd5c0c7ef47906b5f852f2fb099c;
mem[208] = 144'h0968f2baf53704400e2ff927fdd4e1b1f008;
mem[209] = 144'hf8f103e2f57b0a4d07fe0dba0285fc4cf44a;
mem[210] = 144'h0ef407b70525073908c00b7df399f400f80e;
mem[211] = 144'h01720185f21ceff9f02ff8860593069907cd;
mem[212] = 144'h049eed2dfd93fd26049604a1f8c10c83f8cf;
mem[213] = 144'h0bcd0625f5c906a8f2b305a0ffe4fc26f926;
mem[214] = 144'hf3c0070dfd6c0210f7e80f580859f369f90d;
mem[215] = 144'h06f60791f8a50cd6ef73fbf3fc6ffe9afa39;
mem[216] = 144'hfa1e0704f461f9860e41fbac098302eff5e3;
mem[217] = 144'hf87cf4b3fa34fa5a0298fccaf1500f6aff74;
mem[218] = 144'h00bafd21e7f3eb83db9bebaef8d602bc03c2;
mem[219] = 144'hf108f95605540b20fd490b14fc8a0079f4c5;
mem[220] = 144'h0ea1f11df6dfeaaa003bf91beffc0ceffd04;
mem[221] = 144'h03a9f4e202f30d8203bef44deffffe50fa90;
mem[222] = 144'hf3b005f6efbdf937f87f01790c3fff45fb7c;
mem[223] = 144'hf6dbff000772f6d801b4f218efc2ec14f6f8;
mem[224] = 144'h01fb042efc0205bcff9205a8f7f6e923ef65;
mem[225] = 144'h049a071a08e6f4d004d2f40e04daf0060a68;
mem[226] = 144'h0d74f9c50b7af723f9950d9ef1cef070fd4d;
mem[227] = 144'h01cbf4bde3adeb6afc7a0d8a0475f5a4fc4b;
mem[228] = 144'h0b90f781f9def38af77ff35a0709020df3ff;
mem[229] = 144'h0254f708fe0c019bf0a7f06906e00245f574;
mem[230] = 144'h0adafd13f7ba0bd80f180d66f842f2e4fde9;
mem[231] = 144'h0c6408960e26071706c40edf05f407d5faaa;
mem[232] = 144'hfe2f06d60aedf96cff8e0bc0f3ec05b0f772;
mem[233] = 144'h0dd1f6f5040f0ee1fa7605520c22f406062a;
mem[234] = 144'h04f0e489e780ef3febd0fdf1fbf3f322025c;
mem[235] = 144'h0564072eee45015c0667088afbc4fd1efd1d;
mem[236] = 144'hf0160aed05360458ffda033cf218f445f824;
mem[237] = 144'h06470f90f77f09a60026f03e084ffd3bf695;
mem[238] = 144'hfa4a0483ecc6e9060180f9f9ebf6e60de68b;
mem[239] = 144'hfde701e1fa7e0003038dff0cedc5e9a3fe37;
mem[240] = 144'hf21d024d0ec5fa0dfb1ffe9e0e25ffbaf589;
mem[241] = 144'hf8560c7a03810b5cfacb07f30a95ffecf144;
mem[242] = 144'hf1a3099f019803130bec0e62fde8f483fbb3;
mem[243] = 144'h0e48f5a50d22f21507540305f148f2e5f7f0;
mem[244] = 144'h0f7501ddef620b290a3f0c3ff7450623004c;
mem[245] = 144'hfa03ef9804890210085bf369fc430483fe10;
mem[246] = 144'hfe240b67fb9f0d1a016efcfafb490458efcd;
mem[247] = 144'h0488f77c02eaf1f20624fa62fe1ef3e80450;
mem[248] = 144'hf619029a0dc8facefe7d0367f6a60e3ef1bb;
mem[249] = 144'hf979f93bf56f0ac1fcc00333faa20f38f847;
mem[250] = 144'hef5af1b4ff7ff7e705f5eff7f814f851f27a;
mem[251] = 144'h05f80d13f64a00f9fdc8f23701d10a42f846;
mem[252] = 144'h07e2053af8d5efcb030ff17fffc1efd6f0f4;
mem[253] = 144'h07b4014800a4074605daf6b40f72f97b08fa;
mem[254] = 144'hf2f5f6b708ce07e2f9a5071703a90835fc11;
mem[255] = 144'h0f21f66efa57f847fa420cbe02b6ff3701d2;
mem[256] = 144'hf8700622fc6af6570f29fff20a16026cfdb2;
mem[257] = 144'hf586086b091c02d9f19b0459ffc30b910068;
mem[258] = 144'h0cddf98f0d20f58ffbfcf21bf90006c6f1c8;
mem[259] = 144'hffd8f71eefcc01e7f0930da4fef0f54b0a8e;
mem[260] = 144'h0ef1ff20f881f0cef4c10271030b0213efc1;
mem[261] = 144'hf909fa8308e205d605d00e2e0c8e0d17f40f;
mem[262] = 144'hf30a04a3f4b8f932fdf807caf887f69afe2b;
mem[263] = 144'h00ce0633fe29f447022702770dbbf7fa0df9;
mem[264] = 144'hfb70f32a045b0769fdf505f5fda9f9200b6e;
mem[265] = 144'h093605b20653f9ae02660f8ff67f0922f198;
mem[266] = 144'h091af882ef3b0232012c023af764085aeb3d;
mem[267] = 144'hfc510d6c0dd303960a72ffdef272fa8b0126;
mem[268] = 144'h0cebfa49f90ff5c2f3d907c50e38fa46019e;
mem[269] = 144'hfe24f08600cffb1efda70c6d006a00120cb3;
mem[270] = 144'h0f94f11efff40d100345f93809bc07cc00d7;
mem[271] = 144'hf6500979f1b3f2da0557024b0f05f83104f8;
mem[272] = 144'hf57509b3f1ae00930fbef1dff053fbe807e7;
mem[273] = 144'hfbc9f6970acdf648fd71f9cff9d20d03f76c;
mem[274] = 144'hf614f8c501d00268098b0e45f65e08d40f72;
mem[275] = 144'h0e18f6c50eed014f0d63f13a0fc5ffb103ff;
mem[276] = 144'hff3008f1f8ab012e05a308fa0b600f30f4fc;
mem[277] = 144'h001c042d06b2fcb103c5f82df3d900250e3a;
mem[278] = 144'h0e24029502ca02d10cbffe0bffb1f7cb01c0;
mem[279] = 144'hf605fa7c09c90bba09dcf4cc08b8007e07f5;
mem[280] = 144'h07e5017afd06f3770f790e8af170f8b90219;
mem[281] = 144'hf74b0a0fff2dfbbefb48fbcaf2a2032e0dd9;
mem[282] = 144'hf1920833007904bffe7af442f71df5e8f098;
mem[283] = 144'h0067feaa05350d3afba2031ff84ffe03ff6c;
mem[284] = 144'hf254fd9c008f04e4fb3300f5084bf8b1f40d;
mem[285] = 144'hfe4d0a42f8490b5900e1065c0231f0380edb;
mem[286] = 144'h0c99faacfb56095bf7c4f2c00047fb1f0aa1;
mem[287] = 144'hff45f949f55a0b69fdce03b8f543009c0698;
mem[288] = 144'h011507240017f6a10badf251efa9f9f3f6a8;
mem[289] = 144'h012cf15905f70978feadf392f524f82e0ba5;
mem[290] = 144'h0fbff8a50b71feae0a22ffe3002003e80231;
mem[291] = 144'hf655fc2cee8ae1aff9d7ee62f917ec2bec70;
mem[292] = 144'hfdf3072cf84f0135f492018cf2c4f16e0090;
mem[293] = 144'h0a50fa1d06fef3dcff0b0dad09dcfb49f8ed;
mem[294] = 144'h0ec2f0ef0152fd0affd20b1dfe6bf555f74a;
mem[295] = 144'hf82b0da2fd6efa2af118045af014fb7e018c;
mem[296] = 144'hfa240ba4f12e0477f95df68402d3087bee31;
mem[297] = 144'h0a7ff96e0972f5edfc7b0b01fe15ff69f46d;
mem[298] = 144'h0952f991e801fed1ed2705ce0199f92fe512;
mem[299] = 144'hff7cf97bf5d4f085efeffea1efaefcb20ad2;
mem[300] = 144'h050dfedbeedbe1b500b30103026cf5aedf6c;
mem[301] = 144'hf71cf1a9091c01dcfc2b080df2c1f9550b5a;
mem[302] = 144'hfbb40a35ee11edb6f865091f0beef313de3d;
mem[303] = 144'hf893f0e900e9f256ffa1fff50376093bf66b;
mem[304] = 144'hf551ef89fb6804ae05ccfacff801fb10f144;
mem[305] = 144'h0d9df4dbf28c0917010d0e73f12df3b8ffd2;
mem[306] = 144'hfa6b0868fe7a0c3f0ff7f22bf080faa6fe20;
mem[307] = 144'h00effb3203ecf327e8bdee5800e0fa4bf665;
mem[308] = 144'hf11f0abef42409e20317f54ffd76f283fead;
mem[309] = 144'h0dc7ffd40aaa028fef7300100381f1cff0f3;
mem[310] = 144'hf8c203dff46a01e50d33fe3c0d230c9f0273;
mem[311] = 144'h01970034f6d80852fa3d038b0d76f3ca0ebf;
mem[312] = 144'h0f24f7c0f2610c2104e60700f23dfc21fcdb;
mem[313] = 144'h0f1ef516f32202e3efd60937fd0406120568;
mem[314] = 144'hef7df661fb7feca6fdb9e921fe95ff47fd10;
mem[315] = 144'hf0aaf2fcf339fb580c6b0ca9058affa0f6c1;
mem[316] = 144'hfccffafdf810027aeae1fc5304aa00d1f594;
mem[317] = 144'h062a08d206630af4f1a5f6e6f9fdf132f703;
mem[318] = 144'hf07d051fffcafdd0ffe3073c05a6f27005ba;
mem[319] = 144'h045bf7a70ce6f35002b5fc1b0833f65e03f2;
mem[320] = 144'hfd23fbadf722f3c80069faa9f8f9f76bf6f1;
mem[321] = 144'h07ee06c609b8f2c40a3209cdf680ee87f18e;
mem[322] = 144'hf72ffa21f519f031f16ff4e90a3203e10d8f;
mem[323] = 144'hf15eebd3fa28ee44fbefed16f371e662e39f;
mem[324] = 144'hf7cdfd2701350415f573f10d0494fbabff89;
mem[325] = 144'h0a470dd8f6510680ff1cfd26fcd5fc620d98;
mem[326] = 144'h0ae8fc260e8607d50d5706d80929fd7e03ce;
mem[327] = 144'hfa75f7affb000c12fd17fad4f2d9f2780062;
mem[328] = 144'h0e68faab0cb30895f909f52e0145fcfbfc1e;
mem[329] = 144'hf7840a610427ff40052af5180fa2f1b1006b;
mem[330] = 144'hfce0e383ecdff9e2022afc9af101018d07d6;
mem[331] = 144'hf9edf08304e1f2d6fdb1ee9106230202039b;
mem[332] = 144'hefe3e808fa90fdeff0930a1b0e250226fdc3;
mem[333] = 144'h0a9cfa1efe610ade0fd10a3005b803d60512;
mem[334] = 144'hf9a40696f128f7bafdd6f95df42fff69e7e8;
mem[335] = 144'h0c7809420867faa7fdbdf118fd1aefe3084f;
mem[336] = 144'h0722069cfdf701e1068c0f77f82ff5900638;
mem[337] = 144'hf4acf403f423f5730fbff496fb50f9d40b1a;
mem[338] = 144'h0e09fb4ff77dfba9f782f93cf5d5f0840512;
mem[339] = 144'h0961073bf84df02cfeac09c2fdfd02c1f778;
mem[340] = 144'h0bf3ee7cf87cf949fdf70a31f4d60ab20ad0;
mem[341] = 144'h00710537f44500070d77f7a0f2580753f65b;
mem[342] = 144'h0c04f68e06f6028ef36b050003adfd88fac5;
mem[343] = 144'hf52af32a029bff150ae3f0aafc4cf241065d;
mem[344] = 144'h0acaf6e00ab6f3c507fffdd603bb028af906;
mem[345] = 144'h0e78febdf188f5210cb9fb1bf44404a30dff;
mem[346] = 144'hf339028fedacfc67fa2300acead3f28cf14f;
mem[347] = 144'hfb1a0adb038902390c35f345f8bf07380c91;
mem[348] = 144'h033cf236f92af25d09db0cde0d32eda10521;
mem[349] = 144'h024a05a7021efbc103ef0c8c00d5f240f562;
mem[350] = 144'hfc7def39f02af93507910d4ef94ffccc047e;
mem[351] = 144'h09bdf9dbff3bf2daffa4f877f4550530fb5c;
mem[352] = 144'h0e8e046defdef486fba9080dfdb6fbcfe8ee;
mem[353] = 144'hf017f7100239033cfc39fc92022400c0f103;
mem[354] = 144'h09f2059d0393f535fdc9f566fd9e0b66fe74;
mem[355] = 144'hf55cf095e8b2f966ff15fea0f16cf50f0337;
mem[356] = 144'h05c90c62f29f07c20569f4af098bf61d00e9;
mem[357] = 144'h00750aaef9250445092d0b9ef05dfc3cf079;
mem[358] = 144'h0400fecff368fd1c079cf227ff77f60af304;
mem[359] = 144'h0d2d08da040dfeb10479075ff21f0dd9f769;
mem[360] = 144'h02d6fd5108efff3cf0a6facc0091f2b0f9ff;
mem[361] = 144'hf5e008690981f1740fc4f3320ae30fc0fc6e;
mem[362] = 144'hf196e9b3ed980220fc1aeac5fc81f42b10aa;
mem[363] = 144'h0dd90113f9700b14f96ef45d04b7f074f931;
mem[364] = 144'hf6f4ff5b080feb69fa60feb0f90ff347fa47;
mem[365] = 144'h0cb1f296f53c05fbfb1bf028f4e7f4ef0044;
mem[366] = 144'h0bd4f98302f9fd80f49c0317f15af0d00365;
mem[367] = 144'h0f7ff3bdf88d0026f0d6031ffe180137ed4e;
mem[368] = 144'h085b033e07c106f7fcc304affcb0f7c8fab4;
mem[369] = 144'hf40bfe710259fa5af600fec702310a62f470;
mem[370] = 144'h0d91f10efde1f2700b1b0782076ef319fb50;
mem[371] = 144'h01dcfc78fed6f3cf02790806f0f7f4d30ca2;
mem[372] = 144'hf9070c45f31cff3ffb4ff1db026400f702dd;
mem[373] = 144'h00c7fd4c0d1a06befc7afc73fba802ddf265;
mem[374] = 144'hfebe05d2f2b90d0f052603a2f99e0d9f0776;
mem[375] = 144'h0ac40cb2f74805e3fc97fbb60731fa2b0aa1;
mem[376] = 144'hf36f055cf04202eff359054cf21dfd00fd96;
mem[377] = 144'h07a00c33fb00fc39f7500df9fa3bfa500ad2;
mem[378] = 144'hfc0906b80d5d063ef1f40afe0f11fb680722;
mem[379] = 144'hf8a902fbf618059b053704ce0241fca8f95c;
mem[380] = 144'hf5f3ffcf07ff067103810034f6e5073f0fca;
mem[381] = 144'hfadc0065fd4d0c9c0976f3d3fed1f41ff90f;
mem[382] = 144'h00310020f8cbf37af48305300224f270079d;
mem[383] = 144'h069203e90044f4bdfe4e0edffb50ff480542;
mem[384] = 144'hf28ff12bfa91fae7f6de0c3ff45f068bfc05;
mem[385] = 144'h0d57fedbf068f87c0fad078c08e90569f6db;
mem[386] = 144'h06fbf4cb036d0cd6fc5d0c2600d90e43fdac;
mem[387] = 144'h09ec0c3403110cfb019900fdff8bf765fbee;
mem[388] = 144'hfdb4f4690444f3fcf98102ae0f150213f0f6;
mem[389] = 144'h03fafea6fbb5044009c5f2e4f086f244fda8;
mem[390] = 144'h0628f898009bf50b086cf7870cc309470636;
mem[391] = 144'h058900aef087f94cfc09fdd90e39f125031b;
mem[392] = 144'hf5ff0d69ff2700dd07a30f280bd2f71e0773;
mem[393] = 144'hf6a203150693f04d0bc5f2260044f27ef2d0;
mem[394] = 144'hfe2bf130fffcf5130987074d047af845f227;
mem[395] = 144'hf8f10e6200edfde0f02403930c86f9be04d3;
mem[396] = 144'hf102fc5fff60fdbdfc3908d3feb8f2c1f1b1;
mem[397] = 144'hff0c039ffe960b8bfff2fb7ef6fcfcfa06b9;
mem[398] = 144'hfa38ff9bfa5bf5b1f9df0a2502b2f314fd58;
mem[399] = 144'hf6dc041d0872fecef7e9f83afde0fbcb0348;
mem[400] = 144'h0d1aee23fed1e8160bb6005f0a9ae266dd95;
mem[401] = 144'h0574f2b70dc9093805890bda027b0bae07f1;
mem[402] = 144'h0c04fd5df782fdaef3ed0b2af83dfb15f504;
mem[403] = 144'h0d280505f9c9fd16fa9cee76f6fa03e7e5a5;
mem[404] = 144'hfa8901bef3cdfb7a04ddfdb30b3bf7fef2b7;
mem[405] = 144'hf810f2b6fe78fe960ab4f9c8fdfef1710144;
mem[406] = 144'hf9f205d1f99bf433f3df0101051cf56afb1d;
mem[407] = 144'hfeb8fe11048c0459052ef3ea050afbcdfe72;
mem[408] = 144'hff74f444ff38f7b3f84d04d2f978f3ebf8bb;
mem[409] = 144'h053f098cf54d057605ebfb4cfa04073cf933;
mem[410] = 144'hed6ff56b12760963f489eb880241ffe401a6;
mem[411] = 144'hfb21fa9fff8ff7c90389f1cdf06001d50bc2;
mem[412] = 144'h03350af3ea6f028de899f2d7f6ad07c4fc6f;
mem[413] = 144'hf634ff700fd40739fa3a0c86fd8401c20ccd;
mem[414] = 144'h0622fe9cec8fed3d0670f2b7eebb03440297;
mem[415] = 144'hf65a0b0ceef7f102f241fc29fd42f479f221;
mem[416] = 144'h0d16eed3e83de4040999fbf2f5f9e540ebc5;
mem[417] = 144'hf387000002f803590d4a0ec0f2f1071ff7d2;
mem[418] = 144'h0b50f60b0d4c013b0d3f05330791f26dfd6e;
mem[419] = 144'h02fdecdff68eebb1fd89feaff054ee37e45d;
mem[420] = 144'hfdddee8cebcaec2905dbfd0c06a4f97cf5c4;
mem[421] = 144'hff70f0b9f9cdefcb063c07abf37b0e99f261;
mem[422] = 144'h005e0d93fe6001e60eacf5c406def6d107d9;
mem[423] = 144'hf1a6058000a80ac3f0e70cdffdfc0dddfbe5;
mem[424] = 144'hf20609280263f014fc3ff3450d010b8ded61;
mem[425] = 144'h00920a500cad02b6f1e80954f02bf90cf800;
mem[426] = 144'hf012fe22edaaf823ebdfe79deb3109f9fd66;
mem[427] = 144'hf5fcf118f73bf70108e9ffbdfd84f94ef264;
mem[428] = 144'h05bbef5507eef55ef612070006a30107fac8;
mem[429] = 144'h056707ba08c00cdd0b0e060cf97108360082;
mem[430] = 144'hfcfb07a7ebe5fce50655f2f30922f335fc2c;
mem[431] = 144'h07b2f7ffff3c04fff686000afa26f545fd63;
mem[432] = 144'h036204210959002d0e450c470aa3f91901c1;
mem[433] = 144'h0ebaf26b055f05e80455071d047af547f0bc;
mem[434] = 144'hfb7008510681f2c9f5d5098d0e89f9f90e93;
mem[435] = 144'hf63df6ca048cff8ef105f52b06340c6a0728;
mem[436] = 144'hf4d40b5a046cf8ec00e90d000c0cf90a0729;
mem[437] = 144'hfa7bff19f8e3f04afa230a740ae60488fe3e;
mem[438] = 144'hfb0bfe65f3420a2a05650f70f693094f0695;
mem[439] = 144'hf17f0ea8f29f09b003d8fa4ef4f0f7ccf5e2;
mem[440] = 144'h0db005d6f9d6f85af285fea80d0d0244f7c8;
mem[441] = 144'h097f09b7fbdeffe9f167f268075bfee7f978;
mem[442] = 144'h06820a3ffc78f8e30362f958fb6e00e00328;
mem[443] = 144'h0b1f0967f192f5f5f7d7f9cf0ee3f9270bd1;
mem[444] = 144'hf986ff48ff3405affd78f2b5fbf8f10c0f1f;
mem[445] = 144'hf87b067ef95c0cd90849f624f3e1f13ff247;
mem[446] = 144'h0fd80daef397fcaef19df2b704fa0136f453;
mem[447] = 144'h0175071efbd50b14f9c1089cf39d073a080f;
mem[448] = 144'h0e5ef4cf06c7efdaf2fff7ddefbdf2b2f8ec;
mem[449] = 144'hf3b2f51afd6b05e9046c03a4f1c00d840987;
mem[450] = 144'hf42d045e057c02cb02d4f317f2960ad1f44f;
mem[451] = 144'hf1470aa9f7f1fbfef25407d9f801f10df574;
mem[452] = 144'hfc2fff4409c9fba0f41ef418f83ff401ff02;
mem[453] = 144'hf7400b5c053a00df033cf1400ca80247ffb6;
mem[454] = 144'h018df7a20e58fba50b6a061309c7ff7501cb;
mem[455] = 144'hf843037f0e2406bc0323f08ef107ee2109e6;
mem[456] = 144'h0b5c05960218044bfbd8f0180ccdf75ffe3d;
mem[457] = 144'hfcbb05050bef01df0b84f8a1f3aa0df9f5da;
mem[458] = 144'hf9e8072e019004fff63ff7e1edd906240162;
mem[459] = 144'h0b28f5210216f4e9fad2f6340613f8db0505;
mem[460] = 144'hfc76ff99fcdaf496068bffd1fab8fb98f13b;
mem[461] = 144'hf84bf5ddf57d051a05c3f8e604610627fe75;
mem[462] = 144'hf63fee520469fcdd0b39068c0be3079d06bc;
mem[463] = 144'h0a68fe61ee900db60bc8fe19f38809ddf751;
mem[464] = 144'hf9b6ef84f0e8016ef1bbf538fad6ed68fcef;
mem[465] = 144'hffa407c106620dc4fc2a0aeefb4ffaabfb6e;
mem[466] = 144'h09c10ac4fc8dfd0c09fb00b4f07a082a07c4;
mem[467] = 144'hfa7500e7ec60edf408c309fb0785fbf3ede9;
mem[468] = 144'h0bbcf7b9f18df148fbd2094305f0f68b05a8;
mem[469] = 144'hfaeefc450596fbe9f32ff9adf5450a4f0a24;
mem[470] = 144'h06c1090e084fff72f1aaf94b05e0fa06f9f7;
mem[471] = 144'hf4daf0e109a905be059d0d99fe3e042ef12e;
mem[472] = 144'h05dffac9fbd4007ef544fb8df6dcf251031e;
mem[473] = 144'h0eb0014ef814059f0e5406b8f3e9efe900b2;
mem[474] = 144'hf89f0884f625f57df076f4b808bfff42f98d;
mem[475] = 144'h018defe6043af58cfa5c0be1003b04870c7a;
mem[476] = 144'hf03700db000e0414f027f8c1f4b20891f8d1;
mem[477] = 144'hfd9dffcef5810bd7fc970bb206690779041e;
mem[478] = 144'hfadefed0fd940c95f6d50b070ceffa7df169;
mem[479] = 144'hfa8a0cc8056c0a12f926fab60bf70b0ef027;
mem[480] = 144'h0cc70f48fcdff8c4f5390513f18af539fe95;
mem[481] = 144'hfb8bfaabff08f3cef0d7fc15f917031b0918;
mem[482] = 144'h05c9f6a604b8039af85bf1defd76f62c0ac8;
mem[483] = 144'h0f20f847f218fc34ef9b07a0f4f30c7805f3;
mem[484] = 144'hf26ff2eefa92fc0203140562fe2cff23ff79;
mem[485] = 144'h0f5ef9b5fec60d140a660a3e070ff85af73f;
mem[486] = 144'hfb84fd550c4cf837ffa30570070df21901c2;
mem[487] = 144'h04ab08f0f1d003320f3b04d1fcb9f869081f;
mem[488] = 144'hfa200a440412f9f3fa26fa7af65b05caf874;
mem[489] = 144'hfe59ff3df703f0b60e9903440d890077042c;
mem[490] = 144'hf24b03e900320820f0d507c60d9ff5e400c9;
mem[491] = 144'h0ac9090ef51dfc1cf180f6a7fd6c03a0fcc8;
mem[492] = 144'h0068fc4cf9dd0f380f7c04e4f4f3f9aa09a8;
mem[493] = 144'hfaa3f22903320def0289fa39f605f98dfc7a;
mem[494] = 144'h0e28f605f2f6efed04d2f9c8f00301f0f1dd;
mem[495] = 144'hfe070c59fdc6f11406570a08f6b3fe94009a;
mem[496] = 144'hf000f6970ea205e300ddf82efa080b5bf961;
mem[497] = 144'hff09f9c3fd15036b02f90cc207b707660c26;
mem[498] = 144'hfdcdfe06fe60f14a0f8b0a09f20ef5900d10;
mem[499] = 144'hf8f5f3bb0f72fb0c03ce065ff0c5f434055b;
mem[500] = 144'hfbe6f1aff6a4084a09c30d6607ac052e094c;
mem[501] = 144'h0819f7ccfb7ef39b022c00a4f1c50546fb77;
mem[502] = 144'hf568038c057ff6c3ff9d025e07de07b1f6e7;
mem[503] = 144'hf61c031d0eaf049f016dfddf0c9b0219f023;
mem[504] = 144'hf96903eff7b90b1afc620daa00150eb0fa70;
mem[505] = 144'h064bfa00fd85f6eef40a0f9800790cd30efe;
mem[506] = 144'h0ec2f8daf4dd0b4c03bcf35407780e47f43a;
mem[507] = 144'h016c06ab01190e90f49af2320d7df434f3c6;
mem[508] = 144'h04a20b40f9fef1cbf8aafc09fc6af29b0d7c;
mem[509] = 144'hf71ef8ae0ac5005e0bd8083d04990d81073e;
mem[510] = 144'h03a7ff8b023defb505fdf9fdf2d605990525;
mem[511] = 144'h07c5f54f0c630106f4c80a3504fd07f4efd7;
mem[512] = 144'hff5d0f1ffd3f0c10f210f50b0c050366f701;
mem[513] = 144'hf1e00a310f9cff9407580924f2090bca057a;
mem[514] = 144'h0e4e076d0fadf188fe1efb0ff3ff0c94042e;
mem[515] = 144'hf6a904daf698f46f0a1affc4066f0430fbb9;
mem[516] = 144'hf0ff0e00f27d0d56f29101c90074efe1f518;
mem[517] = 144'hfdea0d790ab2014ef8780783ff26f0cafd39;
mem[518] = 144'h04c8f5b40a45027e027b0a2700ca0e6ef4d3;
mem[519] = 144'h08efff000619fc18fa7107e70133080ef257;
mem[520] = 144'h03100a690843fc560860f9f50089f08ef2f5;
mem[521] = 144'hf1b3ff6602eef43e07580740f4b70cd7f4c3;
mem[522] = 144'h02c2fb52f84eee880c3c0d5dfc04fc51f551;
mem[523] = 144'hff4a02410ed0f737f88d04ebf97b0590f3aa;
mem[524] = 144'h0a70ef46f672001af42afdeef6a9f53b05d1;
mem[525] = 144'h0fdd0fdf0978f5bcf9e2f669fe1a02de031b;
mem[526] = 144'h0530f08b04aef612fcf7f771f436ee240282;
mem[527] = 144'hfdf60aa601ae0492f221f96b0af80248039e;
mem[528] = 144'hf380fb82efb8e9b2eedef8c40081f4ade1a7;
mem[529] = 144'hfa740f22ff7200b704c90cd60759f907007c;
mem[530] = 144'h0e3ef329f2adfe5df7090a76f23a07660197;
mem[531] = 144'hf26afadfe6cbffc9ec8d02a8f631f23ef47a;
mem[532] = 144'h07b2ed48f48c0a55048af38ff822083109ed;
mem[533] = 144'h09abf8d5f433f658f024fb88f0d9eda60a4e;
mem[534] = 144'hfaa2f751f6ce09a70cccf7e9f0b4f020007d;
mem[535] = 144'hf731f74af66602af0382f1adf780f433f2f5;
mem[536] = 144'hf805f113fcacf4e1fa410267eef502a70446;
mem[537] = 144'h0031fd96f58205210ee406550c07f0b60c6d;
mem[538] = 144'h0351e9a9fe66f2f9fdddf209f8e80057ff49;
mem[539] = 144'h0416fc31f7fafeacf228061ef8cefedbfd28;
mem[540] = 144'hfd03fdc9ea1fe7810277e8a207efeb3ef578;
mem[541] = 144'h0a4c0ee60b7c063e03370ce0f350f37f080d;
mem[542] = 144'hfe570123073ff83cef92fc5a061ce148f3cb;
mem[543] = 144'hfdca08bc0a20024b00b00aaff6aefbe0f4f0;
mem[544] = 144'hf9b1f62b0124f99ff2b4f98cf368f4d2efb8;
mem[545] = 144'hf86c0ecaf3a4f6faf1a1fd1df72efd930a81;
mem[546] = 144'hf0cffe0bfee80a35f5e60726f6c107c106b0;
mem[547] = 144'h0b27f0d602fb00210377f60ffc8c0327076a;
mem[548] = 144'h07ee022df372f74c09a9f6e5ef95fc5802bd;
mem[549] = 144'hfebb0927f80cf2b6f512f6b6029a0969f5f3;
mem[550] = 144'h00990b9e08b1fcf307a3f762feb5f5f2f8eb;
mem[551] = 144'hfea5ff130016f22e0659f6e7ff220c680bd1;
mem[552] = 144'hf944ef39f91af11804b30668f00209dcfdba;
mem[553] = 144'h043901d8f1d4fca5fb2c04a5fca1fee70da0;
mem[554] = 144'h0260fd4bfcaef27ffa010a880221f128fb72;
mem[555] = 144'h08cf057ff069f23c0b19f92afc6e0da40399;
mem[556] = 144'h01590441fdf00298fd64fea80a64055feeee;
mem[557] = 144'hfc10f0990b7708b60c49fad9076afc43f1c4;
mem[558] = 144'hfd90eecdee5007ed09c2fbab095c0436018e;
mem[559] = 144'hf1b0fd29fdea02650702f0ddfcb4004cf38b;
mem[560] = 144'hf418f95cfd05f4130001f02df80ef676fca8;
mem[561] = 144'hf7d202400b580785f4b3f1eef699f3daf130;
mem[562] = 144'hf8b4ffa3062906530651fac6f679f666f87b;
mem[563] = 144'hfc50eeeeee51ee44eae9e9dcf572ee4607bf;
mem[564] = 144'h094ff6fbfe6fff8a06ae01defdaef7adf4bb;
mem[565] = 144'h00bb0c3401bb0af4f179f3bcf40c0a59f8b8;
mem[566] = 144'h03cef3f3f7befff20c18f87e05f7f49d02f2;
mem[567] = 144'hf855080e0e3ef69bfc1a080ff6e6fcdc077f;
mem[568] = 144'hf8e8ef91f2f3f2670be1f5c7079c0608ffcd;
mem[569] = 144'hf979f83004e7f39bfffb0271f91ff4180f58;
mem[570] = 144'h056eede0ef59ec97f6d8e11ef0f1fbb80cde;
mem[571] = 144'h095a07eaf5f6fb3af168f7dfefd0085bf931;
mem[572] = 144'hf86a080bfc63ee2b03c4007d09f3030b0659;
mem[573] = 144'hfecb01bd0a7cf3730e8503c3f574ff41ff37;
mem[574] = 144'hfcf9f1effab3e70e030cf533fee0fdd5fe47;
mem[575] = 144'hef4f0a2601f30897f75d06ac0949f75fefd3;
mem[576] = 144'h029504b905a6ed29f180f74cf7b9f0b8f6ea;
mem[577] = 144'h0e47f74cfab8f81a07e30ce3f036fe73f228;
mem[578] = 144'hf21c06280e2101990bfef6b5031cf599efa7;
mem[579] = 144'h015204ab0470019d08daf951fb08f732f6cf;
mem[580] = 144'h0444001b0ab90bc10cd2fbceff95068ff7ef;
mem[581] = 144'h0745f9d1f4dcf2aaf57cf8d9f1940eab05fa;
mem[582] = 144'h0599f8c207600513f56cf6d2097bf652febe;
mem[583] = 144'h0882fb030ee6f9ce0ca3f744f4e1f0e00090;
mem[584] = 144'h0c66093a037bf7c2f2bcfbf7fe5b0d5700ee;
mem[585] = 144'hffcbf344085905b9f9b9f6e9fbe503fdff63;
mem[586] = 144'h0acafc99f268e902fa23ef2bf37b07e106df;
mem[587] = 144'hfd7bf4e2fc330a170770fd8af6bb098c0af7;
mem[588] = 144'h04bd0296fe7e0036081900e2083006f7fbd3;
mem[589] = 144'hf09d0de4043bf0aa0c920e64f6640e77096d;
mem[590] = 144'hf313f9c60ae50890f67d06e5f6f0f10ded75;
mem[591] = 144'h053c0a0ff21407fa096afe090b6dfef8013f;
mem[592] = 144'h04ecf75bffddf1ee04fb05710c860c660669;
mem[593] = 144'hf0f3f933fa01f619ffaf034ff3f9fe42f0bc;
mem[594] = 144'h0a5b0db00428f66c089bfad5fc5a042af82e;
mem[595] = 144'heff2ef9e05deee94fb57f1da0a470503f4a3;
mem[596] = 144'h0e430a0605ce03a1fc50fb4dfffff6e1f2a2;
mem[597] = 144'hf862f7d3fdc808a7f458f8f9015c0bcc0178;
mem[598] = 144'h0d6ef725fc4707baf1e80f13fe83f9a101da;
mem[599] = 144'h0ab60cd308790bfcf2b60b26f9e1fc3a08cb;
mem[600] = 144'h0d01f292fdc809d2fef8f359054c0d0b04f4;
mem[601] = 144'h0b8e0e9304220403f395f564f9ab0c10ffae;
mem[602] = 144'hf8db08aa093004f50a13f935f431ff8c0426;
mem[603] = 144'h05bf0029f732ef87f16f0e12f5affcccfa82;
mem[604] = 144'hf265057df164f9000dacf341098c0b0d0d52;
mem[605] = 144'hfa1604d0097efd34f950fd8d078ef540fcc8;
mem[606] = 144'h01250b4feeccf2a8f6a109520bda0d1a0200;
mem[607] = 144'hf547f8b2fcde0dbd0473083f010bf324032c;
mem[608] = 144'hfb22f35b07a7f248026d0f69f219fcabf9dc;
mem[609] = 144'h0cff058ffc140be3fc4c0802f6b1f416fa5a;
mem[610] = 144'hfcaef4f603bf046af85dfeb20741f38f0112;
mem[611] = 144'hff3df7ffefd90ca2001903310c02fc4df345;
mem[612] = 144'h030f09440b84f5b90c33f0eafff9079705ac;
mem[613] = 144'hfc5400c807c3facff8ddfd63f491f3f709a6;
mem[614] = 144'hf2c6f884f05b008ef89c0e35f29d0b86f485;
mem[615] = 144'hf9aa04e9f198f67ff136f5ba034f0b9a020a;
mem[616] = 144'h008bfab3f117052a09f5f4210314f548007f;
mem[617] = 144'hfd1af237042e08e80a2af17d092808920c47;
mem[618] = 144'h069cfd9d0710f11c064dfbd204330987035f;
mem[619] = 144'hf9a6f568f782f31cf2700d9ef6460d85f4a9;
mem[620] = 144'h06140ac90bb4f272049e0e4b0c20f8e0099b;
mem[621] = 144'hf17d0885061c03b500dbf2c006e4ff0fff6c;
mem[622] = 144'h0be5f79f0838f1fd0d2f00f1048bfa53f336;
mem[623] = 144'hfe1ff19cf0d8f68fff5006ac09e50833f9ea;
mem[624] = 144'hf1a2015707240bf7f244f830090cf710eed8;
mem[625] = 144'hfbc0023d0b87f077f8b8024cf6ac040ef424;
mem[626] = 144'h026ff169046bf1720f8900d50e6affc4f61f;
mem[627] = 144'h0a2d0e2d0906efd9ee1bfab3f741f756fd60;
mem[628] = 144'h0bb106ac0a300a05feb9084afd17f8630cbc;
mem[629] = 144'h07c902a308d5f24704d8f0e5fb7af478016b;
mem[630] = 144'h004af052f4ae03a7f6660c7a05b4001dfebb;
mem[631] = 144'hfcf900c10088f81df84af94bfed1f1130c2d;
mem[632] = 144'hff45fc4bff820d25f1360554007c0653f435;
mem[633] = 144'hff550fb5fee30c8a075703850792f37d05f1;
mem[634] = 144'hf993f532f0bdeeb20837043df48dfabceb70;
mem[635] = 144'hef97ef8808d30cf2f84bf36af8adf7f80cc9;
mem[636] = 144'hfa6c0149f5d5f66cfdc907c4f41402790ddd;
mem[637] = 144'h0a1bf2b40de50666f876f816f581f7810fb2;
mem[638] = 144'h09fd0c430d5109a8f190f0adf98b0eb306a8;
mem[639] = 144'h090cf14c05ca0ef302a406ed05f50448f0f7;
mem[640] = 144'hf17af60afd320ee4f79703c4f57607f50375;
mem[641] = 144'h052af64200e3f116f5d00fc80ce40c5d0fd2;
mem[642] = 144'hfaf60371f4d90710f168fcce07f005b60d2e;
mem[643] = 144'hf19ef01a0b3af4e6f5f201f005f90b3f0944;
mem[644] = 144'hf1730184f0130ee6f0cff76c0481f1550210;
mem[645] = 144'hffac0181055cfafef33dfd9df62709660adf;
mem[646] = 144'h030ff336f53df365fa6ff1130a3a02b3fcbe;
mem[647] = 144'h0dd4028d02490a67fa3b0fba08c6f1220a82;
mem[648] = 144'h0c020f83ef750e1203ec06900e6d0243fb96;
mem[649] = 144'h09820de908bb04be02deff9dfea6f19af3a1;
mem[650] = 144'hf8c9f0ce0d3d05d40742024af852ff1efeba;
mem[651] = 144'hf01c0dad09e5f8d4f6e5fa9707070dbc0e81;
mem[652] = 144'hff62020e08d00e67f6f0f9820ca8f8f90916;
mem[653] = 144'hfa320993f05d0ee80ae20819f643f578f810;
mem[654] = 144'hfec50bb508dff816091bf7eefeddf136f810;
mem[655] = 144'h0746f5af051bf92802a10a8bfd220100070f;
mem[656] = 144'hf193f71f04faf694f91a0f140410f0b9eb27;
mem[657] = 144'h0e7a0e7ef0cafdcf0e31f51bf854fc64fca2;
mem[658] = 144'h0efdf7b3f7c6fd7cfaf8080cf226f456f31f;
mem[659] = 144'hf952059f0842f8ec0298fb6bf600fb7efb47;
mem[660] = 144'hef8af93bf7fef65b09e502af04acffbc08d0;
mem[661] = 144'h047df284fa670a2afd11f045ee11fd79fd35;
mem[662] = 144'h07920435feb1f69e04cef9840dbe01dbfe06;
mem[663] = 144'hf67002ef077dfe0e0772fcbc09c9f92d09d9;
mem[664] = 144'h03820ef0ef46fd2209effb6afbacf913f3b8;
mem[665] = 144'hf19e0151f173fc6d024102d20967f8f00662;
mem[666] = 144'hf4e6f404fab3ece3f43ff791f323f55bfad0;
mem[667] = 144'h0dc7f44301d70e57fadcfb66f8c30caff260;
mem[668] = 144'h05060054fbdbff78f04cf13cfbd0fbbe0460;
mem[669] = 144'h01dcfc34f4d80685032a09a30b1503370b96;
mem[670] = 144'h003704a907e1f24107300841f85de997ff4c;
mem[671] = 144'h04560b9c094a0ced030909e2f0a602b80ba1;
mem[672] = 144'hf22f0e16fd98f90af401ffbff715feed015e;
mem[673] = 144'hf2fdfabaf7e6f20cfca506a6f302f56907ad;
mem[674] = 144'h034f01dd019a00810589f0db0bacfb99f81f;
mem[675] = 144'hfbf307460aebf101f16e0659fdaa0488f7a6;
mem[676] = 144'hf6140ae0f074f6e9013407d404e8fb830379;
mem[677] = 144'h0c89011fff7cfa40f1810deb099508b907f6;
mem[678] = 144'hf57f0618fbe8ff49ff4cfaf8f379feba05db;
mem[679] = 144'h0898047f0a840e5d0caa0e0bf8d5fd9ef56c;
mem[680] = 144'hf485f69d026affc40a2cf0040978ff0cf063;
mem[681] = 144'h00720b27f0e5fbf6f8100c7c007d0ad109fa;
mem[682] = 144'h0999f40f0b52f023f1adfb6500e80544fccc;
mem[683] = 144'hf38e0e95f3b0fdad003d062cf671f8fd0ed4;
mem[684] = 144'h002c04eff66df7260d16f515f721f1290edd;
mem[685] = 144'h0094f1af00fefce60b2fffaf0c6803e40507;
mem[686] = 144'hfe82f3b4ed49fb49fafb08befb5fef8604c7;
mem[687] = 144'h0dd401c20a07017d003cf0f6f334f2a3008e;
mem[688] = 144'hf076f9930e5701b407a9f9a2f67007ba0b0b;
mem[689] = 144'h05eef4ca07280f57f473f555090cf96f062f;
mem[690] = 144'h055d05b6f7b80d29f1d0fbfdfb9b09ddff57;
mem[691] = 144'h073ef2a60b6cf773fde301d4f30af0cbfbcb;
mem[692] = 144'h027807d90582022cf917074fffc80a330f17;
mem[693] = 144'hfab0ff17f9960dcf01180e320ce503730fce;
mem[694] = 144'h01af0fbbf6ae041bf6c5f6da0dd5f23cf7db;
mem[695] = 144'h0423f42204dc02e307c00fa00509fd6204af;
mem[696] = 144'hf38efbc506b6f1d3fb42fb1c0feb0a92f735;
mem[697] = 144'h03cd0342f123f6fbf20d0be4f1fb060005aa;
mem[698] = 144'h007f0c010d1d074100910156f24e0243efba;
mem[699] = 144'hf824fff600490d72ffb6f213f6370ecef352;
mem[700] = 144'hf877fab4fa51f81402970bbbffc503f1fd6a;
mem[701] = 144'h0edf09600e500ea8fc50fa5df82c06cf0db7;
mem[702] = 144'hf6360f76fc200237f49c0ca4083f05c9043f;
mem[703] = 144'hf49f0bf303f2fc5e0a300acffce9f42902dc;
mem[704] = 144'h0f280e470971090ffe42031bf6ea0a91f221;
mem[705] = 144'hfd32fa82fdd6041f0152f289055cf1df089b;
mem[706] = 144'h0ba0feed002107fcf1bff5f909810d17051d;
mem[707] = 144'h0ed506b50a2d0b960424fd88f972045af44c;
mem[708] = 144'h08abf21df6fa06d8fc690a0af313f15603c3;
mem[709] = 144'hf96ff8940ede079001490246fe13085200ed;
mem[710] = 144'h06290bb3f4600bbf0a980f7e075bf658f767;
mem[711] = 144'hf7eff902fcb5016f00d1f948f3e6fe8af22a;
mem[712] = 144'hf4b2f620f7700bb3f52902590400f704f77f;
mem[713] = 144'h040afdcdf413fbc0fdf30d940c1e0dfcf801;
mem[714] = 144'hfd5af188f343f35afdfdfdc40751fee4f1a2;
mem[715] = 144'h0bdd0e21f5a70bc2f82cf12803ec0cd10483;
mem[716] = 144'h00eff6cf0647ff6204a2f26600910d10f04f;
mem[717] = 144'hff21f4b0f821f8df048cfff70c4f0ea5fc34;
mem[718] = 144'h0b8af25a05260cf6f24cf9fdf12000670c5d;
mem[719] = 144'h0613fe09fb21ffb7f093f216f07f08d30a61;
mem[720] = 144'h0783fd07f3fe0987f08e01630f3ffc5202b7;
mem[721] = 144'hf393f39ef85d0500f0f8044a039af1df0d2e;
mem[722] = 144'hfd71051109a30ec90213fbe7092af5160aa7;
mem[723] = 144'h0f00f1250bbbff1bfcf5fa2b0ec8f156fa8e;
mem[724] = 144'h0be3f0f9feba03b8f9c3079d09d40bc6097a;
mem[725] = 144'h03c60f3bfdb304180a6108a2fba80dbbfe61;
mem[726] = 144'hf0c0f13705faf576f707f9cbf9befcb3f400;
mem[727] = 144'hfc680b39fc0b05780ebc0ccf083bf6090c64;
mem[728] = 144'h0ed1f5b1086cfa16010400dcf7fd0e6bf556;
mem[729] = 144'h0113f1db0190fb8d019bfcc3f85df95d0b5c;
mem[730] = 144'hfd15fee504620b1ef38609e4f3d4f1890ab2;
mem[731] = 144'hfd3908f3fff1fd180db9f251fb84f656009e;
mem[732] = 144'h043afb040a2801d906390d24f7f80751f676;
mem[733] = 144'hf2a3068e03ba076ffdf0fcf6f83e038a020b;
mem[734] = 144'hf08ef75ff37608ab08b1f1bb0cc509ac06de;
mem[735] = 144'h08b1096a0355f5a10f070e67f91d0b58fe07;
mem[736] = 144'h07fff01af7640b7405c2f427fbd4f2ae026a;
mem[737] = 144'hffb80891f5fdfa670171019ffaecf0a1f9cb;
mem[738] = 144'hf25609d30537083b04d2fa93fa9007690433;
mem[739] = 144'h03cef15a013f0a86f027f1b2fcc906b1f743;
mem[740] = 144'hf2540ab8f14bf09208eb046dfc24f1fa0ba0;
mem[741] = 144'hf5b9f667f8a90ccefe91f94dfb40049b0af3;
mem[742] = 144'h0688064104f90646071d0681011d01b8016a;
mem[743] = 144'hf832f5f6f19ffaadf7da0aa9f0a6f11105e9;
mem[744] = 144'hff79037cf754ff7207f5f7100baf03f709f6;
mem[745] = 144'h0ca0f9e106f1fbe20495f315f7c3f004f97f;
mem[746] = 144'h09d506bb0df1f585f641f9e507c0fe96fd19;
mem[747] = 144'h083f053a072f080afd6cf58c06c507d8efbb;
mem[748] = 144'h06f4f257f86606c904e90211055007be0cc9;
mem[749] = 144'hf91a0e47ff000d0bf485019bfdfaf7200ce8;
mem[750] = 144'hfae80f630e0200e70fb1fc22f62c0ee50528;
mem[751] = 144'hf2dcf9bf0dbaf5b2ffddfc30052df42f0518;
mem[752] = 144'hf110f9ecf41609850c2701ab041ef87a00a9;
mem[753] = 144'hfec5095cf6ddff37fcb008b60617019df68d;
mem[754] = 144'h0be20b67f12dfe04f795f0970e6601c809d1;
mem[755] = 144'h0b3f09370c2800b30609fe2d0d810f57fc07;
mem[756] = 144'h0b3202c70ae4f977f02ef32bfbe70ac20e9c;
mem[757] = 144'hf6c8f7fe05a4fab204f4f2fcf935078e078f;
mem[758] = 144'hfc14f332f73c019f052bfe790609fdc90187;
mem[759] = 144'h0cb1fa22fcd30f7a0214054dfec7041bf66f;
mem[760] = 144'h042a0e2f055f0344f8ea0f5df1cd026e0343;
mem[761] = 144'hfc28f023f39307fefdd506baf00b06cd0b85;
mem[762] = 144'h0700fbb4f307f8d4035101300a3a02b8fed6;
mem[763] = 144'hf8c9fa0cfa4efd89fc4e0945fcf6fda60c2c;
mem[764] = 144'hf5fcf3f7fee8f7ee0f720a3af1bd0d38f69a;
mem[765] = 144'hf56e030a08ad0a44020df6770cd4f8abf505;
mem[766] = 144'hf874035b0946f2c9f75905400f3b08befdab;
mem[767] = 144'hf4acf0cc00eb0baef2ec066201c004eff71a;
mem[768] = 144'hf3c0f4dc009fefe5f476f4c5f15408b4fdef;
mem[769] = 144'h0c1002c9ffd2f0840854f1bdf77301faf23c;
mem[770] = 144'h063906bef6a4fe92040e05ec0a64f5d301ed;
mem[771] = 144'hf8f707f9f48c07b8f47cf5a703c10570f4a4;
mem[772] = 144'h0d83044e01dbf2df06da0fe4f9db05b9f98d;
mem[773] = 144'h09970dc0fde9fb990ea90bcd0a84f755fac7;
mem[774] = 144'h0ea809d3fb0d0db7f72d0e1cfc31fecaf2ea;
mem[775] = 144'hfcbb08d7f68efcec031b04f9f7d60915035a;
mem[776] = 144'hfc95f4f6f3f5026109ccf797f632fd5b058d;
mem[777] = 144'hfbc308130ca8fc37fd2d0dc9064cf9760f96;
mem[778] = 144'h02990070f9380afb04d20c060de9089def16;
mem[779] = 144'hf4fdfaec09b0f54106cbf24f0dabf8aef33d;
mem[780] = 144'hf2d50b76f1070d3bf7af096efdf0f9e50370;
mem[781] = 144'h02f8013208f7002c072f035b010ffe37f90f;
mem[782] = 144'hf4a8f929fc3307680562f7a2f26b069a0700;
mem[783] = 144'hfb25f2d7f7cc0395fa23fba8fb09ffd4f8b7;
mem[784] = 144'hf8540fc1f1a60c9f09daf846f74a0ddb0dda;
mem[785] = 144'h051cf283f106f65ff52ef170f9cbf9ad02a0;
mem[786] = 144'h0aecf868fce1005c00f6058304180607ff94;
mem[787] = 144'hfbd20f290881f654f4ae0628062d0756fd39;
mem[788] = 144'h00f7028df87df3c102cdfd48fcc402f102c1;
mem[789] = 144'hf34e078f07b0058906a3fb1f0ef2f2bf0d77;
mem[790] = 144'h034cf22b07a802b3079cfc2007cd0d44fa28;
mem[791] = 144'h0bde00f809ac0e8a05c7f7dd070801bbf055;
mem[792] = 144'h09380ae800a0f9810794febf0d7c02dd0095;
mem[793] = 144'hf3a10e6c0f23f49ef17af593fd37fd30fd55;
mem[794] = 144'hf9a8f98cf61cfbbff0150cb1f839ef4cf47b;
mem[795] = 144'hf903fa8004930bedfac1fb6f0f37efcbfa44;
mem[796] = 144'h09ba0a42fa83f538f22b08d00abd09090b36;
mem[797] = 144'hf4540a8c00c2f954f758f1400866f180014e;
mem[798] = 144'h0e61f2f6fbd2098706390df9f6d7f14ffbb3;
mem[799] = 144'hfeb4f9aefe710f680727fbd0effaefcfef8c;
mem[800] = 144'h0be2f758f42fec82f71f00e8072af24aec11;
mem[801] = 144'hf8e5f614fbe30b58fee10292fb0707020078;
mem[802] = 144'h0590f9600d49f77600710aa0f8c3f7c606f0;
mem[803] = 144'hf5b9069ceda7e543e4fcfca4ff7df5c6e199;
mem[804] = 144'hef09f31f0c0505c203e1f1c1fe51fd41f7ed;
mem[805] = 144'h043dfda4f6edf64b038504a3f59c06bc0466;
mem[806] = 144'hfd6c0452f3090dec0c670c740e1dfe75f4ed;
mem[807] = 144'hf362fb2af4df08c702e6f3790a82050907fc;
mem[808] = 144'h05db0575f2df053ffd8b03bafc92f50df917;
mem[809] = 144'h0e550ee90740f25cf4de02950a32f9f80e37;
mem[810] = 144'hf007ea44f5abf157fab9f32d02b0fd510a3f;
mem[811] = 144'hf7c5faf70314fa07fac9f867f3a2ff89f8f9;
mem[812] = 144'hf8faebe6fbbcf9c3f95f0875faf5f717ee9c;
mem[813] = 144'hfb6e0c4cf400fb92f16a020ff432f4ec004c;
mem[814] = 144'hf980eb70f19cf78af39afcc2f27f04d5e798;
mem[815] = 144'h0a50f23f056ff3bb06e3003304ba000df1d7;
mem[816] = 144'h0edd00f50ebef085f0b80a07fe220c26ffb1;
mem[817] = 144'h04f808c3fb5df21502dc084af6af052a0434;
mem[818] = 144'h066ff5f20374fe110673fdf5037803e8fdd0;
mem[819] = 144'h0e9904f4008e0083fe71f712fb3e0ba0f3f1;
mem[820] = 144'h0b4e03e4f0aafcec09f20787f84af660f10e;
mem[821] = 144'hf581fd010642f83af0cafb64049104fff032;
mem[822] = 144'hfb7f049909d80be60702f7cb0bc7f6ad0ae8;
mem[823] = 144'h05270cf5fc310e55f9ac0e7ff1a8f651eefa;
mem[824] = 144'h0685fbe5ff76083cff8e0f9908490a34fe8f;
mem[825] = 144'h0d750a24f33d06b008bd0e4cf4a900e50bb7;
mem[826] = 144'hf10ceed4ecdcec5ceed2f07e0c3f0140032c;
mem[827] = 144'hf30cf4510dc00b66009df8a3fdb30ab4f2b0;
mem[828] = 144'h02a900f1fa08056af62d091a07a30086f10e;
mem[829] = 144'h0086fb9bf94b0adef8030e360ddcf23904dc;
mem[830] = 144'h0ab40226f6c1f5d90aa8023cfbb3003af992;
mem[831] = 144'h06f1fc26ffc00efc05270f3009110651ff32;
mem[832] = 144'h0fa0f7e6059b068400f006feee31018e03ad;
mem[833] = 144'h049bfb3df8c5f9ecf2a1f5d305820de10302;
mem[834] = 144'h0ca4032ef6fcf49dfbf504570f67f728f158;
mem[835] = 144'hef9b0ccb0dbaf1bc0159ef09fc83ef6bfb44;
mem[836] = 144'hf4690b93f08d001bf2140fd2fe380588f3b0;
mem[837] = 144'hfb74f91805b405bf029ff53afd6305610c4c;
mem[838] = 144'hf11d0640fc3ffba4fcfcf3120fd0f875fb19;
mem[839] = 144'hff80f20af871fffafa560990051bf1cb0a5e;
mem[840] = 144'hf38df81cffb60f37f4d40aa6f7d2f999f9ad;
mem[841] = 144'hfe65f28c0517007bf4770433f1f7000efd55;
mem[842] = 144'hf36ef80eef8c05c70525f34a03d40479fbc0;
mem[843] = 144'hf99ef53bf077feef0d9af81d06d7f6120c70;
mem[844] = 144'hf216fbd70343f4540b2dfff8f0c6fe1b0016;
mem[845] = 144'h0ee5f2c0fde5f78ff176fe2700120d690163;
mem[846] = 144'h04dff18202af02c8efb1ff0a04f50bf503c3;
mem[847] = 144'hf8eb0970fe4508dffd3ef898f021fe130651;
mem[848] = 144'hfb100c230ba400ec0db3fffdfea90f54f07e;
mem[849] = 144'h0cb00ab2f8380a39ffa000d10779ff62fdfb;
mem[850] = 144'h02a808c2fb0800bd03a40544fad7ff690f5b;
mem[851] = 144'h0568f332f37df7a6f09c08080be50bf7fc55;
mem[852] = 144'h090efbcf0325f7f4055e0147f04c00cbf8f8;
mem[853] = 144'h011106780232ffaffed90361fc94f670f487;
mem[854] = 144'hf58dfefcf95efd9c068ef6bff745f0110084;
mem[855] = 144'hf36e08acf09af37ff4eff8470598fc98f4d2;
mem[856] = 144'h0d7c08a40084fee90decff620f03f96403f4;
mem[857] = 144'hf7acfb640a4807c10c830bbc021307390d88;
mem[858] = 144'h07c80e280c11f636f6ce0ea803d9f6aef8ed;
mem[859] = 144'hfc29fb56fa38f00303f30d07fd40fbfff996;
mem[860] = 144'h01430351f9100c8bf38ef57cf17ffbd00848;
mem[861] = 144'hf73ef18df04302b60591086707dcf4770b3e;
mem[862] = 144'hfaac0f19f2d1f7d6012f0bd3f0baf56d0e06;
mem[863] = 144'h061cfc6ef4f3006af15e0a9efaad0c12f139;
mem[864] = 144'hf85aecebf0c3fbc706e00c9007fafcddf564;
mem[865] = 144'h0c1cf41807bc035f08760223efe7ffb5f3aa;
mem[866] = 144'hfa41f2f6f87cfcebf9cefb4af6ea06c5063a;
mem[867] = 144'hfa82fda2e909dfc1edba0b480402f85bdf1c;
mem[868] = 144'hf7f5f60409db08ccf9840299f2b50837ffe5;
mem[869] = 144'hf6ab0a9af5c90d2ff4d4f22109990b4dfc06;
mem[870] = 144'hfcaef3150a6df6a80dc9fecaf47b09acf9d8;
mem[871] = 144'h051ff7b8025201b903000003f042f855048d;
mem[872] = 144'hf9f8f8b107f4ffe7f289f5fa01ec051e0a98;
mem[873] = 144'h0020f818082c00ad0269f062fb0ef8d9f165;
mem[874] = 144'heba3e770f645069ff28df0f5fdddf758fa37;
mem[875] = 144'h062dfdc3f265f996032a05c6f34e024806b2;
mem[876] = 144'h0c4b0549f180ebc7065ef49dfd0b0862030f;
mem[877] = 144'h0622fec1fa7f082f0b99fdb2f6dffb74f19b;
mem[878] = 144'hf079019ff938e683eded0b16035a058ae4c7;
mem[879] = 144'h0096ff15f04cf7cf0af8f08eeea2f0e1edc7;
mem[880] = 144'hf5e109e3f8f5ff95fcd00e6b0b43f3a309da;
mem[881] = 144'hfab2063af41d0d05f4280314fb2e08f60842;
mem[882] = 144'h0fc6fd14fc50f1bff2f9fa2cefec03cf0281;
mem[883] = 144'h064bfaccee16f6a9fa960195f2f6f873f206;
mem[884] = 144'h0471f415f2cef3a106a2f4a4f314f2a7f493;
mem[885] = 144'h06cbfd9bf1d7fa630b770e3bff7bfd71fa63;
mem[886] = 144'hf7990948020dff900da409dafc330d530c33;
mem[887] = 144'hf2320b87f76c04770278f1abfe81f7cefb72;
mem[888] = 144'h0ee3fbd6088b05790cb9f0d6fd14f78c0360;
mem[889] = 144'h0c0cf4c10da104160c08f24607c204a6069a;
mem[890] = 144'h0a630163ffd8fb180000fa20027f05def030;
mem[891] = 144'hf8330389fa530436045ef882074ff0f4f0b3;
mem[892] = 144'hfd1df5e2024d0063ef07f64b0a7df79af906;
mem[893] = 144'hfcb0f0f8fcfe03dbf117029ef58f0c940fdf;
mem[894] = 144'h0011f8ef0375f742f5d5f8e5ff4aff9507f0;
mem[895] = 144'h0135052cfe5e0ba8fd79ffb40bb3f619f36d;
mem[896] = 144'h0797fd78f5b0f1f406d5fecbf8ddfff5fc46;
mem[897] = 144'hfda3f60f09aa0c46065ef149f79102350f4a;
mem[898] = 144'hf69f04280c05fba00536060f0d0af7d8fa42;
mem[899] = 144'hf358ffeafef50bb2f366f9ddfadf09a1037a;
mem[900] = 144'h0b9604d4faf0ef97f3170448fff30aa300f2;
mem[901] = 144'hf9e30817f63602b1f42f03d4f6c500e4fe63;
mem[902] = 144'hf40609eefb150a4502130480f266ffd5f393;
mem[903] = 144'h06fdfaac04e0048e09e7fd3cf3cdf3f3018c;
mem[904] = 144'h00600e1e02acf1e3f312024a0dbbf3a7031c;
mem[905] = 144'hfd42057b0e7308ecf18207a40cf001a1fbf0;
mem[906] = 144'hf3adfdda036f057dfe5b04520c96fb90f406;
mem[907] = 144'h0f100b6ff091fb3ffe02f3800b42f55ef2b8;
mem[908] = 144'hfcb4f94c0d4af2bfffbf0f8efde6f494fa3b;
mem[909] = 144'hfe5f0c9df86c0f1a0955f2bc06b3051b0441;
mem[910] = 144'h0360fff10a9c064e0c82fe130e9e0bba03a8;
mem[911] = 144'h0dc50aadf15ffbe0f27e0a4c09deef400082;
mem[912] = 144'h06f80ca10d4df74cff55f933f75501d9fc63;
mem[913] = 144'h09b8fcb2f9baf7d30a91f89a0dac0879f47c;
mem[914] = 144'hf928087c01c1f327f0eaf0d7041404c802b9;
mem[915] = 144'hf2580d030169fdfd0b0e0deb0ac7ef12ff96;
mem[916] = 144'hf47c001bf7e602580647014c0d970e5b047d;
mem[917] = 144'hf12501850aee0b8cfe21f8dd06830377efd8;
mem[918] = 144'hfdbb0441009ff52ef10a01dc006405060ac1;
mem[919] = 144'h01930d65f12e098af6f0f8e4fe6201720e1e;
mem[920] = 144'h0057fde80d7af34c0852f74efba0022606d8;
mem[921] = 144'h06e2f15bf6bff3f8fedf0a2ef2b8ff4ff411;
mem[922] = 144'hfafbfffb0a38ee34eecdfe65f38eecddf919;
mem[923] = 144'hfee1f610f776f5afff98f7b40b54f4dff505;
mem[924] = 144'h0867f7590ee2f3acff5f0c840d8bffbd053c;
mem[925] = 144'hff34ff56f220f6fe0ef9f5590d6a0409fd3f;
mem[926] = 144'h054908e40b78f6150cd0fb2d0db80763ef37;
mem[927] = 144'hfb6c0a87f343f1040ef800caf0f0093b07fc;
mem[928] = 144'hf5fb00be07e6f360fdfe0da10a790b79f18f;
mem[929] = 144'h0d7ffac3fad40e880036f59a08590d4d0a26;
mem[930] = 144'h0a990070fa5f0382fc4b0e0a090bfa590c7c;
mem[931] = 144'h01b00c06f3a7f6480afe0abbf850f62ef43a;
mem[932] = 144'h0b820983f3230343efeaf8c6fb18fb5dffec;
mem[933] = 144'h09c0f307f5a9ffd20da3ffdafd8a0581f3ea;
mem[934] = 144'h0f8ffa32f9d60cd2f1c805b9f243f980f870;
mem[935] = 144'h0f7efbd7f5290a32f581f8bc0cc0f9d90381;
mem[936] = 144'hf378ff84049afd09fefefd730267f3d201f1;
mem[937] = 144'hfddff10e05d702b6f346f8a8fe8df891f90a;
mem[938] = 144'hef6b0296f6bbee080900ffb1f44907130c39;
mem[939] = 144'hfc320ad70260ff58f8e604a802c8fe210d91;
mem[940] = 144'h09e80b2f082f041c0aca0aa9f48b097df7c5;
mem[941] = 144'h05e8fdbbf1fb0f8f0b4e01a3f1980e93037a;
mem[942] = 144'hf2bb0b3204a5fbe8f147f2bef955f2d30a18;
mem[943] = 144'hf2befc26f03df0b6f7980c8608310d20efbf;
mem[944] = 144'hfde00bce0e5d0f9a0e17ffe1fdd4023c0230;
mem[945] = 144'h0bba0d7e0512fe75f01e00ccfc18f6a80c22;
mem[946] = 144'h08a5f17f04c0f726f24e040c07f5f3cd0af2;
mem[947] = 144'h0c8ef6caf27bf9f7fd34fd9ffdcefebcf93c;
mem[948] = 144'h0b6c0006fbdcff4afcc405050dddf5df0be3;
mem[949] = 144'hf16cfcbbf0b4f3b502d3065ffd23f1e7087c;
mem[950] = 144'h0184000eff990b38f5f3fa6e0d05f48cf7a2;
mem[951] = 144'hf1e80d730105f5a8053c0d93f087f9a3f1c5;
mem[952] = 144'h0479f1d8f2c1f9ea0e3bf26cf5a8009e0c05;
mem[953] = 144'h04b2f2710d8c05420ca7f527080107880669;
mem[954] = 144'h0b9bf827f906fa9efa73f1070bdf0bc10af8;
mem[955] = 144'hfb9e051a036c0b69f3d9010e0a6ff30df5d7;
mem[956] = 144'h01180d2c00df0ebefa2d0063ff77f0a00982;
mem[957] = 144'hf9c30824f6bdfc320ee3f39c07b602370fea;
mem[958] = 144'hf57af8c9fd66ff41f9100ca7f648fc3b0314;
mem[959] = 144'hf9cff142f35dfc220d8cf9200da7f2650c04;
mem[960] = 144'hf167fb1c054df22f02820c12ffcd0ead0b8d;
mem[961] = 144'hfff60abdf13f0c5dfb62077205c3031af22f;
mem[962] = 144'hf664fe150382028ef956f45103a404a90bbf;
mem[963] = 144'h0336f20d0d55fe79f34ef3bef9a10b640212;
mem[964] = 144'h07a5f50df95a0f310a470f1ef919fe49f238;
mem[965] = 144'hf938f9d90a25095af71a09230d290e29000f;
mem[966] = 144'h0025f415fe0ff2adfbeafe78ffe3f6f4fabd;
mem[967] = 144'hfef1fbd103770237f9f5f8540cfb0466f5d7;
mem[968] = 144'hfa89f9ccf1e60b60fd2f0bda02f3009003e8;
mem[969] = 144'hfb6ff6d3f56903060e62f2daf43109fdfae4;
mem[970] = 144'hefc3f57703a10ea3f73d080af64bee580a02;
mem[971] = 144'hf3d203f60d38fe2efb960800faef03290219;
mem[972] = 144'h0922f920fbacf2710b7cef91f1d8fd290456;
mem[973] = 144'hfba300970dc40e97f87b082a09f8f919042f;
mem[974] = 144'h0fc20c0cfd86fd90fb540149f6a8f190f86a;
mem[975] = 144'hff8ff68305b50eac07bef753f4010416f023;
mem[976] = 144'h04f2fcaaf58cf12008caf6c3f5e1f40af606;
mem[977] = 144'h02ac041c0889fec60eeb0d0d0659fed3fedd;
mem[978] = 144'h086908e7f2b7fa8ff6d20e03f5bc0de8f28b;
mem[979] = 144'h097df68d0c0107edfe7403adf3c006e8002a;
mem[980] = 144'h053108950a5dff3009780021f711fdd5f00e;
mem[981] = 144'hf992f7f7f2d9fcc807a10043f494f1d00582;
mem[982] = 144'hf98ffcb508f40d4f01b70545f48d01adf4f8;
mem[983] = 144'hf162f6a4011ef2fc06a207ebf9c7fcaff182;
mem[984] = 144'h0f42f3b4089dff7bf5bffeb30194f849f7e2;
mem[985] = 144'hf44605d7fd53fe5b09830edaf2d8f892f3a9;
mem[986] = 144'h0916fd65f0f80c0c07dcf5320b0bf12bf882;
mem[987] = 144'hfc8efd1e01e2faf1fda9fad205e40de00a48;
mem[988] = 144'h0ff2fde9f20706f8f4b0f16e033bf77d0386;
mem[989] = 144'hff1e0c0ff35500b9f90a0cb0f71cf4ceff96;
mem[990] = 144'h02460072fddeef770e460efb0f53f42d086d;
mem[991] = 144'h0a7e005e01ddf586041c0e1ff0fef2c6007c;
mem[992] = 144'h08c9027bf774021c06caf3a9f453f6caee2f;
mem[993] = 144'h0d7d0b8e060a02aef47bf0e602ac03410771;
mem[994] = 144'h03a30f9cfba407de0714fee90a2d094707fc;
mem[995] = 144'hf04d02b903b8f0d904baf361034207b501bc;
mem[996] = 144'h0c73095806f8facdf995f63ff21bf174030d;
mem[997] = 144'h0026fc2905fdfc1c0c65f28aef56f58503ab;
mem[998] = 144'h020802a300d20e510531fa58020a06e8089a;
mem[999] = 144'h0ee70312f1d40975f43e04230a2dfd89edb4;
mem[1000] = 144'h0f08ef65faf60218046d011501a3fee4ee95;
mem[1001] = 144'h00710b1d0841fe74fa4cf11209a1ffb8f2ee;
mem[1002] = 144'hf7e4f7c2f31ffd7df3c4007a08d2e4bc094d;
mem[1003] = 144'h0a750d0cf6ee04350d38f71cf22209a8000f;
mem[1004] = 144'h0eeffe060487f789f2e7ef5c0ef8076efd28;
mem[1005] = 144'hff5bf068fe8c08bd027bf5b005cc0f14f1f1;
mem[1006] = 144'h0f1d069df9b80966071b072bf026edc0fc7b;
mem[1007] = 144'hfff608fffeb3025f0653042bfa26016cf209;
mem[1008] = 144'h0b8e0cf8f17efa4bf47cf3fa0c7afd9af35d;
mem[1009] = 144'hf54ff6eb0dabf05908c50a5e0e8ef6680748;
mem[1010] = 144'h0ed40b280e0d08f8068e0dd806c8f49afce4;
mem[1011] = 144'h031cfcacf0ea00a0003cf9070577fb4ceff0;
mem[1012] = 144'hfc0f01400291ffea0434041602b70c3cf3a0;
mem[1013] = 144'hf36101d4065cf324fc360551fcfbfd8e07cf;
mem[1014] = 144'hf9fb0bd1fd420e350cf1fbcef315f566f21a;
mem[1015] = 144'hfde4f733f31afa0bffe1fab9f209f2f200a0;
mem[1016] = 144'h0e1af3f5f754f57009a3f38cfad9f6e90c6b;
mem[1017] = 144'hfc54f60603bbf4d0f87e0c2f0968efe305a6;
mem[1018] = 144'hf040055af9a7090c0417f5ecef68f8e8f216;
mem[1019] = 144'h0e32000def9bfe56f2fd041ffa74fc78fab3;
mem[1020] = 144'hff670120efeb0afdf39bfee6f29807cffc3e;
mem[1021] = 144'h0f310ad0f82ff7e005fefe7ef46204d70aa6;
mem[1022] = 144'hf76d017bf93c0ca1fc94f317fc440153fe43;
mem[1023] = 144'hfe6f06fd0d2305de0cbb0753efd3f81d004a;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule