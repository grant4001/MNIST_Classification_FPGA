/*
Copyright 2019, Grant Yu

This program is free software: you can redistribute it and/or modify
it under the terms of the GNU General Public License as published by
the Free Software Foundation, either version 3 of the License, or
(at your option) any later version.

This program is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of
MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
GNU General Public License for more details.

You should have received a copy of the GNU General Public License
along with this program.  If not, see <https://www.gnu.org/licenses/>.
*/

`timescale 1ns/1ns

module wt_fc1_mem7 #(parameter ADDR_WIDTH = 10, DATA_WIDTH = 144, DEPTH = 1024) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'hf799fd65f5bef039097ffbbc099e079cff0b;
mem[1] = 144'hf690f638f196fb84ff5f01c0f6010906f545;
mem[2] = 144'h06bb035efa7af4d50015f6f50bd10d740252;
mem[3] = 144'hf5ebefa1fb8ff5e4f7b7037e009b014c0eb8;
mem[4] = 144'hfdb90107079fff79f5b700700ea50a5d098f;
mem[5] = 144'hfed3f411ffc2f7240a450f21fbadfed707c6;
mem[6] = 144'hfab300650073032304e2f66206720014068a;
mem[7] = 144'hfc3306d6fef4f13004a8f00a0dbe048cf0fe;
mem[8] = 144'hfd3cfa550f47fa6a0915f6f3fd5204ff09d1;
mem[9] = 144'hfb6d0a0cf0650508f7c70dd403bc0bb4069d;
mem[10] = 144'hf24208bcf09d0bc50302095d0cabfe47f390;
mem[11] = 144'h08b400ea064f0a350ac6f71afa7ff898ffa8;
mem[12] = 144'hf75e0ab50cf80e7701480cbc0c88fc020efa;
mem[13] = 144'h02ae06230d3ff667088c0f53f41df2cafb2e;
mem[14] = 144'h0a570a4a0230f911f8ff05daf35cfddbf0be;
mem[15] = 144'h00560141020f0df4f4c4027cf07a0a83f7d7;
mem[16] = 144'hf0c6039df6aefbed000ff4db0c1ff49bf366;
mem[17] = 144'hf30ff98efa16f52ef4e307c3f670f00e0015;
mem[18] = 144'h0f6308bdf0c20915fa69fc39f5020fbc0fb3;
mem[19] = 144'h0df2072c0815f35902f809c4f310f7650371;
mem[20] = 144'hf7c0046bf0b00f620878f86afd440273ffd9;
mem[21] = 144'hff36ff5f09a3f160fa0af5b00a61f82701f4;
mem[22] = 144'h018406580ca7f1a50ce40edbf7bcf9bf08ec;
mem[23] = 144'hf7e3fc86f414f713f90104d8f0640cd3f2cf;
mem[24] = 144'hf98bf6f1f9f1003d03ba0267f7800b9ff130;
mem[25] = 144'h022207c40cb30444f5e50956f0df02e6f708;
mem[26] = 144'hf2050938fddaf3eeff14f717f1910e23f728;
mem[27] = 144'hf5410715ff1f0589f9770dd2fe6609270006;
mem[28] = 144'hffdb0082f09afabe095f09200bbcf6a5f727;
mem[29] = 144'hf1e701730910fdeb00b7fdd101a401f101a6;
mem[30] = 144'hf96ff346f04ef90efa390186fea5fb0700e2;
mem[31] = 144'h0a7d09c302fff3d50b4705fdf860095e009f;
mem[32] = 144'hfb47f71900b60636ed1ee817ed17f0f10c07;
mem[33] = 144'hf0890eadf9a40c68f8eafdf801d1fc0300d1;
mem[34] = 144'h0b97fb0fefcbffb2fd130b760bb50116f15b;
mem[35] = 144'hebe9ff52008d0c86f0b1e743070aec08031b;
mem[36] = 144'h07e1ef3c03ad0d13002d0092091cfe680ad5;
mem[37] = 144'hf9fcf162fd10f841ffaefb2efda400c2f3f1;
mem[38] = 144'hf2020836f6f6062ef63d003dff6002a0fa20;
mem[39] = 144'hf284014af00ff8a9fb6cfbe8fd7f0eaf0850;
mem[40] = 144'h0680ef63f6bbefbdfce7f82f0152fde00e94;
mem[41] = 144'hf652ff28072c029bfe89f930fdfaf641fcec;
mem[42] = 144'h0901015a01d0f812f684072efa0e04f30221;
mem[43] = 144'h075802fbf23e03020c6df76df7eb072b02bb;
mem[44] = 144'hf2adf84b07b4ffe804b20f06021802620dc0;
mem[45] = 144'h09fef794009df52008e7f8baefe4ff480c38;
mem[46] = 144'h039af0e5f1190ac4e513f5f4eb890030fe36;
mem[47] = 144'hf9dc0a13f87e051deb45fad2f64efec2ffc9;
mem[48] = 144'he39deea6f299fd10f96df715ec2c004afdfe;
mem[49] = 144'hf01ef44fff85fd92f31ff2d1f6f8055d03ed;
mem[50] = 144'hfa9df4ee08e4fc52f7dcf21af60600d5f1b2;
mem[51] = 144'heae2f407f19bf315011706070101fd810c54;
mem[52] = 144'hfaea0b960aa4f4430552fb58ffe8f608fea5;
mem[53] = 144'h0eb30ace024cfe1cf017fbc50aa10daf0378;
mem[54] = 144'hf9ff04cbfd9408a1f391041900d8ff9e0dea;
mem[55] = 144'h088ffad8fb2bf07a020bfbabffe9ff58f035;
mem[56] = 144'h091fee75fe1108060813f248ef14fc9b09f2;
mem[57] = 144'hf82801e4f82bf139f59def66fe59fe34f864;
mem[58] = 144'h0fbde94de87bee6df3fceb07e7c7ff70f2c8;
mem[59] = 144'hfe92f586fa5504f6f818057ff211f1ee07cf;
mem[60] = 144'h045f08f2f181f1e400fb0cec0846f813f29e;
mem[61] = 144'h0f67f3980e42f93f0a1800ab03e8f2cff408;
mem[62] = 144'he119e7def77aff25f7c3e835e24cf954fa7a;
mem[63] = 144'hf09907e505830c7cf233ed69fd49fabf0527;
mem[64] = 144'hf396ed2bf708f181f400fa6ded4c06f00510;
mem[65] = 144'hf88907adf150054ffa0bf7520115f11a0ed3;
mem[66] = 144'hf4cafaf9f657f2a703e1eec60449f6210e28;
mem[67] = 144'hf553f01d0af8f8ec01600345f6160731fcef;
mem[68] = 144'h099e06580b450e93fee1f6e1f58ff39b0e0a;
mem[69] = 144'h02e1f3100356f9d9f5a80b3900aaf40e03ac;
mem[70] = 144'h0d06f8c5ff2f0a16039cf579fc7df3d3f08d;
mem[71] = 144'hf2ebf9aff50403d1f179f4a7f7caef07f7ce;
mem[72] = 144'h0552fdd5062a0553f974f5c20796083bf940;
mem[73] = 144'hfc3ff95104ae01e80da7f5aff8c104800d39;
mem[74] = 144'hfc97f46ae87fec0feafef4e80a0ff999045a;
mem[75] = 144'h0427fe080262f999071d03970563f2e50bce;
mem[76] = 144'hf84ff4eef4edf1f4fc71ffe60552f48ff9f4;
mem[77] = 144'hf3de0975f1d6fd41f972f4daf33d0ca2fb36;
mem[78] = 144'hfa3b039f0477fb54f365f844eaaf02c7ee75;
mem[79] = 144'h0442f58bf386fc79fd440565f5b6ee4cfcac;
mem[80] = 144'hec05fc51042b098ff35be8d4ff170a8e0733;
mem[81] = 144'h0182fadff302f6ad05180d360183fde60234;
mem[82] = 144'hfb49f1a6095403c10c96056c03b3092cfcd5;
mem[83] = 144'hf702ee4bf765095bf271014df4ecfa0a03bc;
mem[84] = 144'hf166fab9f91603e8066ff920069205fbf20f;
mem[85] = 144'hf07cfc3200880a03fa69f2250a2301760aec;
mem[86] = 144'h0ad60e6109c20c66f09bf26f051609a5fa7a;
mem[87] = 144'hf22e06510849fb05fae008670b110cd8f77a;
mem[88] = 144'hf759fa28fd3f0868f34d0111f815fc0d0256;
mem[89] = 144'h0aa90a37f2f6f26801cdf553fcbff85c088e;
mem[90] = 144'h0bbdfef8f8e509a6049cf7b7ee9803fff069;
mem[91] = 144'hfbc30da10b6afdc001a5f380f9cff7df07e1;
mem[92] = 144'hfe080acb07e5f2fc00d0f82708d6ff2df08a;
mem[93] = 144'h0196096508530d0df078fa11081af41af56a;
mem[94] = 144'h00b101f1ed4f02ba0585ed3e0464ed8d0aea;
mem[95] = 144'hfe6709d8f841083ff8fc0b51f025048ef41f;
mem[96] = 144'h01360e02f33d0515f2570727fb800687f8ef;
mem[97] = 144'h0a89fefbf78efee20058029dfa76f5840275;
mem[98] = 144'h0baffd90096cf39ff888f8ebf459f70f05d0;
mem[99] = 144'h045903bbfa42f402fcb3fb3e09620940f62f;
mem[100] = 144'h0cf803d9096bf2760cbbfe98031a02f9fbb5;
mem[101] = 144'hf4620551fc82f3f8f0cc0914f018056e0c9d;
mem[102] = 144'hf60cfb510fac05bdfa76fe060d5e0446f964;
mem[103] = 144'hf6290a11ef350197fa8b05aaf368f8fbf5e1;
mem[104] = 144'h08b3f743f446f7d4efb60df3ff13feb2ff8b;
mem[105] = 144'h05610c210dae005cfec9083df49507780eff;
mem[106] = 144'hf3cc0772f28205e3058df96a040302dbffe1;
mem[107] = 144'hf1e609380117fa9f04fc03b00deb09d20574;
mem[108] = 144'hf8edf2d60e570bf4f850fff40392f6790c90;
mem[109] = 144'h0e9bf3bbf7190c300ede06230d64ff6e0f4f;
mem[110] = 144'hf06f095b0b390482fa9f00260e3ef0160d70;
mem[111] = 144'h0c72f3320936f6f00c1df48afdfbef5c0ccb;
mem[112] = 144'hfe6effef032cfdd5fde4e87f0be60be102a2;
mem[113] = 144'h0248f27508aef14308ff006f0ee102620dfb;
mem[114] = 144'h00c704aef5fa00ecfd270e2ef73c003bfc54;
mem[115] = 144'hed3f05bbf795ffd8f35f02b7ec96f14b0132;
mem[116] = 144'hf993ff210056fdb6f254086ef50efed501e2;
mem[117] = 144'hf928fa41050cf12cfbc3fc69fb480437f312;
mem[118] = 144'h08ddf4b2fc800cb80c8bf8aa03a2ff6b067f;
mem[119] = 144'hff5b02190901f56ffab4f0b20c15ee4bf8b1;
mem[120] = 144'hfb4007fc0038f8a50a530b15ef7df44dfc87;
mem[121] = 144'hf17a038df80f0413f59af22eef4efecbf203;
mem[122] = 144'hef64f5b1ffd509fcfcd9f6d30436f203ee78;
mem[123] = 144'hfa1dfb25fe7ff246f55df48f0c48f49c0c63;
mem[124] = 144'hf9bc0b16fd870700fc9efd9cf4cf0014f6f6;
mem[125] = 144'hf4e4f913f5f9095efe2af840042ff5d50ded;
mem[126] = 144'hf5b8ec290073fdd6f848efbd072603540e28;
mem[127] = 144'h0527f1dd0e7ef81d06af090dff80f0c9ef1c;
mem[128] = 144'h07d30d1e0c64010e058f082ef1c8f528fbce;
mem[129] = 144'h0328f1e80bc9ffd502650df1f4b7f615f1f6;
mem[130] = 144'h04190034ffbcf5e2fc83f5dff65a03d10fd4;
mem[131] = 144'h0dab071b0cd70bc8f8f80d6101bc032cf34c;
mem[132] = 144'hf51ffb3a0ddbf9be0843fe50fc050aebf6e3;
mem[133] = 144'h00150814fd880cf801e403e80c760bbbf27c;
mem[134] = 144'hf8ae02def1a70b9cf2b80136f5410c6ffd22;
mem[135] = 144'h0bf604870a330ebafee50bc202b7f799f0b0;
mem[136] = 144'hfd6ef89f0d460a1f0506f227052b01c3f00a;
mem[137] = 144'h0fb008cef98e0f5c078dfc2606d1f3d80308;
mem[138] = 144'h0493fbf00e6d038a03def20ff1baf45d05df;
mem[139] = 144'hf2f50580fcbaf3b5fc4dfb9d0bfbf125f73a;
mem[140] = 144'hf05a02cd0462fe88028af5200733f32af5fc;
mem[141] = 144'hf883019404d7f613f55df2c2f4b40603f9ed;
mem[142] = 144'h04250c1d01c3fe97f28ef6c20329fa70f903;
mem[143] = 144'h0746fe3ff70b0db5004600a400e50c2909b0;
mem[144] = 144'hf927f9d3ff6400d402acfe800f79f639093d;
mem[145] = 144'hf6970b6b03eaf87bf1faf8080b22fc3b0511;
mem[146] = 144'h0eb806ed0b2dff8df99e01440db0fe790ac4;
mem[147] = 144'hf73c01bdfe0a0de3058aff78028e0a61f92d;
mem[148] = 144'heff1f673096afe36f2890e65f1e7f8f60580;
mem[149] = 144'h0c0a0ad6f6f80c8a0e530871f8f5f0520116;
mem[150] = 144'h041eff5a0c5604b50172037af753f1430d21;
mem[151] = 144'hfa22021105ad01e5f3dffc8e041ef1a7f646;
mem[152] = 144'h06e407ddf324f428fb8bf6ea01d9f160fa3e;
mem[153] = 144'h0867efb6ff5bf457053f0e150041f3ad04b1;
mem[154] = 144'hf0e5047d0918f6c0f1ea01470211fdb5072e;
mem[155] = 144'h0c75fd1d03b001f30bd2f7acf4e206f3fd96;
mem[156] = 144'h0a15f9b80af8025708930c7af62cfe3bfd52;
mem[157] = 144'hf7e3f72b0c5c05e3f51afcdd08ca07a9f0dc;
mem[158] = 144'h0e1503890d420d2b094e0bc20bd30481f8a3;
mem[159] = 144'hf0f3faa0fec6fe8afb4df622f97002b8fff9;
mem[160] = 144'h0d45f94bfa0804250114f16105480c39f25a;
mem[161] = 144'hf81bf243faa405e4f7f30d2c09300c3af32e;
mem[162] = 144'hf799f98c03f4fab9fcb302b7011107fff7d4;
mem[163] = 144'h04920dc1001bfea20856f57cf973fa1f015c;
mem[164] = 144'hfb7f0f99f8c0f8b705d3fe550f95fff20551;
mem[165] = 144'hf8e00ab008bbf77cf2c50d63faa5f1e50afa;
mem[166] = 144'h01c1f7dc0cfbfce00b7cf969fc54f94d0460;
mem[167] = 144'hfb95fa5508670477fb7df0edf511031a0ecd;
mem[168] = 144'h0ee7f2d5f73e065203c7f8aff48205c6fb8d;
mem[169] = 144'hf9f90bd30bba01a000d80a75f884ffd40321;
mem[170] = 144'h02a4f96ef1e2f70afc15ef0000ebfa420f91;
mem[171] = 144'h0e43fee008d6000ff239f7bcf911f6f502f7;
mem[172] = 144'hf9bd0024f63df1eef9c8f7ab035d0eef0d6d;
mem[173] = 144'hfa7407b007f2f5f20877f2a70bee05d60867;
mem[174] = 144'h0cb80241004901acff330e1f0c54f6fcf21c;
mem[175] = 144'h093bf5770aeef75dfea00b79f9ac00ebf307;
mem[176] = 144'h08e20bfa085204b0ff180ada03abfeaa0fb3;
mem[177] = 144'h04bf0c34f8a307ed0d0a01ca00b6f00f0379;
mem[178] = 144'hfa170690f6dff69d0bfcffc30e500200fd52;
mem[179] = 144'hf751faee093ef853fb38fee0fb6cfccdf5b1;
mem[180] = 144'hfd6f06400fe9f7920cfaf2160073f356081f;
mem[181] = 144'h021c0566f65e0034f0680d5effa100a0f1b7;
mem[182] = 144'h01f40e05f3f80115fd20fa77fa120234fe23;
mem[183] = 144'h08c2f7270880f038f3c7fc2f0465ff50f396;
mem[184] = 144'h066f06540d1a0dfef51309a7f2400dff0697;
mem[185] = 144'hf81df2060f34f5d5083300c8fd09f092f6eb;
mem[186] = 144'h0931f2d40214fb57f326f681f0b401b4fa85;
mem[187] = 144'hf4e70c5df504fce2f9f20faa00590b9b07c2;
mem[188] = 144'hf8e50e070413f28ff44705c30b9407040ad0;
mem[189] = 144'hf999f1dc0d3d0cd70404f65df490fe34f1ba;
mem[190] = 144'heffe04590a190212f15cfb280821f996f4b1;
mem[191] = 144'h024df818f30bf2600a9ff90fffef005d048b;
mem[192] = 144'hee3608870e4bf622fa53f255f11df5a708b3;
mem[193] = 144'hf9e7fc6df0f6fc7a0c63067ff02e05af09b5;
mem[194] = 144'hf8b10d230f12f34c0e52fe19f66408a8fbca;
mem[195] = 144'h0ac3ef16f374f53c0270f0430c5bfaacf819;
mem[196] = 144'hfc56ff0b06e10e72f487f4780d36f8db08ca;
mem[197] = 144'h0d7effbafa480135f6d20de6f780fb140924;
mem[198] = 144'h0b2aff4df6a8f118fd0aefd80219ffa5fe77;
mem[199] = 144'hfeae013f09e7ffdafd6e0bfe0dae0b2ef763;
mem[200] = 144'hfd5a0accf096fc5af42b0dadfe4004c10ded;
mem[201] = 144'h0d9c0145f6b2f1b3f7bb045bf48cf670ffed;
mem[202] = 144'hff7cf3fff624f1dff343f91d04e80242f5b4;
mem[203] = 144'hf97504130098f1d1f2560c8f0ca20e9f06a6;
mem[204] = 144'h01a50d5b0d8bfd5a0bcc01d1f67cffd507e7;
mem[205] = 144'h0eb0035ff144f410f683f0ebfdf8fd160a12;
mem[206] = 144'hf74607d00446f9640670f1ee03f0f1f90724;
mem[207] = 144'h0368f3b1fd4ffd38f2100bcd06f1070d03b6;
mem[208] = 144'hec1dfa0803b508b5f7eaeb14eb9a06a1efbe;
mem[209] = 144'hfdbffd850b5700d20f050542f764f900f102;
mem[210] = 144'h0c760583ffcaf2d4ed2bf21d01d904b8086e;
mem[211] = 144'hee23f68bf37104cef0500388fd88ffd4f6b2;
mem[212] = 144'hedcafafcf6fb09e80d170107f69903bb028d;
mem[213] = 144'h0b9b0b02fa2b026eef4a0b47f39cff2eefec;
mem[214] = 144'hf27e0bb20076f3860402f1810d73051c0bba;
mem[215] = 144'hf14d0536005af84af2b6fd3c0718f29ff572;
mem[216] = 144'h082bfa4e05fafa81f0f3eb7bfd38f2cbf78e;
mem[217] = 144'h0200001d0db608820c5ef27cf61af89d0ed7;
mem[218] = 144'hf2e6e97df52decd4eaf7fef2fd62f1e0023e;
mem[219] = 144'h014dfccdf62ef0fdfe7907090710fb8c03a6;
mem[220] = 144'h02f90342f4c805f20aca09dcfe4bf32ffb69;
mem[221] = 144'hfbf8fd7a058a005c08aff5a002010c7ff5df;
mem[222] = 144'hf129e6fefc23f39503cdf7a4f6d2f76c0750;
mem[223] = 144'hf9aef316017cfcfef12906910b050506fa35;
mem[224] = 144'hfe7d0acbff70f59101b4ecf4f88e0be10c61;
mem[225] = 144'hf23cfac4f7e8073ffa23f4340fb40a4000b1;
mem[226] = 144'h089df2a909430ae200a8f52d06c50c8df042;
mem[227] = 144'h0623ed75f254f38cf53cfc8404dcf0930113;
mem[228] = 144'hf734f4d500dd0c2a0dce0d4d05920ab30914;
mem[229] = 144'hff6405aefd7e012bfe8efc9e02fd058bf936;
mem[230] = 144'h0bb3f3adffbf0220fa330db3f73afddbfbec;
mem[231] = 144'hf97df474f06104f7f89d0107fe47030403a1;
mem[232] = 144'hf38c0d1bf50bf1a20dc0fd9805edf49c0296;
mem[233] = 144'hf25c08dc045a0739f96805fd0774f3c3efde;
mem[234] = 144'hf8effb6fef8efc8dfe0af7c8f68203fb0558;
mem[235] = 144'hf67cef55070ff41afbe403b1ffc3f6c10242;
mem[236] = 144'h0b70f193f45afbb20d55fa590b91fbc1fdfa;
mem[237] = 144'h077f05de0dd2049203270b84faf201a1fc13;
mem[238] = 144'hfa59f62e0321fa39f96ce44dfa2dfdcb0dbf;
mem[239] = 144'hf9deffea0b8a0bdafa5cf878f3ff0ad10026;
mem[240] = 144'hf270fd1bfdeffce40faaf97af07f090b0b5b;
mem[241] = 144'hfe68f0b60f5f03460f3e0e9f069ef931f984;
mem[242] = 144'h0efb05430a0b06d0088c061dfc2b0813095e;
mem[243] = 144'hf6bef669eecaf44ff117f77a01f1f26b014f;
mem[244] = 144'hf7c708f307a80d77fd870314fe820834f928;
mem[245] = 144'h065e06a10a6a0092f69a081203c0fa26f677;
mem[246] = 144'h06c0f974014e0f96f480f58f01e40d2c0635;
mem[247] = 144'hf0dd072f0005f3aff7a30601ffea0dba0d43;
mem[248] = 144'h05f00176020bf3ca0333fe9c06e7f8f20817;
mem[249] = 144'h0cd4032cf8ba06800bfdf8fc0a4407b0feb4;
mem[250] = 144'h0165fc890c25fdbcf4eaf4a2fe3e0598069f;
mem[251] = 144'h087dfa330b600a3bf7be0ef80402f1550d42;
mem[252] = 144'h09030d90f497fdc8fb9af26bf744f19b06e4;
mem[253] = 144'hf2080c140e1a08d7f5f20add073202cafe51;
mem[254] = 144'h08b00c87045e036c04e8faf7f863eee60571;
mem[255] = 144'hf38ff02c063e0e61f7daf08f0d52f76ff7b7;
mem[256] = 144'h0867fe8df5a1f789f84802fd06570a9b061c;
mem[257] = 144'h0f5d070df3ee02950377fd26f689fc630511;
mem[258] = 144'hf526fbf101bbf00f03ea0e8309c301e4f10c;
mem[259] = 144'h07c2ed770acf05eef4e8fc5af0fcf3ff0347;
mem[260] = 144'h0b13fc7dfe090e3bf79a09aaf7ca098cf806;
mem[261] = 144'h0b97f30b095b0d3f0f0cfc4defb30e870f2d;
mem[262] = 144'hfda7fccef082fb76fe210617f8d40e0df4e7;
mem[263] = 144'hf971fd54006bf066f80dfb47fd5e09b30be5;
mem[264] = 144'hf9b0fbea0b64f2f0f9f9f391f5170d3f0e82;
mem[265] = 144'h04c600510d64f8010a95fc90febe09fe02f7;
mem[266] = 144'h06c9fb82034efd2af72afded071ef34afefe;
mem[267] = 144'hfa88fa5d0162f20ef008f21dfab0fcac0415;
mem[268] = 144'hf396f9760183f9f5fae2075f0d9e0453f84b;
mem[269] = 144'h0ab80f9df3b10845019af4960789ffa700e4;
mem[270] = 144'hff550359fd0107000c4ef5d5035a0b48fc06;
mem[271] = 144'h0e0e01130e4efad1f0b502c2f51d0e980e3d;
mem[272] = 144'hf33dfd8cfe2bf8b5095505a5f6d301260c4d;
mem[273] = 144'hfcc4fb40010bf24204dcf26204830e6b0320;
mem[274] = 144'h09c30014fdb609edf3bd01bcf5360330f095;
mem[275] = 144'h04c0085bf04cfcd309650eaaf1d9fe07f003;
mem[276] = 144'h06eaf34af14af1faf24102050abaff4ef1e7;
mem[277] = 144'h0dbe02c8054cf082035d052f02bc04bdf2f6;
mem[278] = 144'hf68dfcf308310d750f3b05780d5505680d67;
mem[279] = 144'h067c0f7d014c010600cef94f080802ecf405;
mem[280] = 144'hf4df05d20a9b082ff921fba9f98b09cf07b3;
mem[281] = 144'hfec70119f0f4000b0050f15ef927f353ff86;
mem[282] = 144'h0cba0075fd70f083fedbfdd101bcfa14026e;
mem[283] = 144'h0cb5f8fef927f656fecff5360216fa49f720;
mem[284] = 144'h00cbfafa0da1f3640d77f024faec0003007f;
mem[285] = 144'h094ff3f3f2baf0f4feee0406fed1faf6079e;
mem[286] = 144'hf459f1fefa350c9bf599f018fb36f306fded;
mem[287] = 144'hf27df789088f0f71fe31030fffde0586f331;
mem[288] = 144'hfe22fd44ff6aef6cea17fe03ed51f631fea1;
mem[289] = 144'hf07703e2fc03fb40027df2ebf3aa0aaff1f8;
mem[290] = 144'hf9cffb96f8ecf68e04600347f5850242fde8;
mem[291] = 144'hfeab03bbec80f74eeeaa00def7defb60f56d;
mem[292] = 144'hf524086b0de70ccb0a11fff6f844f7160679;
mem[293] = 144'hf792f5e6f758f58afdddf56604250d6e06bc;
mem[294] = 144'hf4a10e98fde3fee40a60fb67f2dfffe3f48e;
mem[295] = 144'h036cfb40fab7fcd5056d0db30b6701b7f120;
mem[296] = 144'h04bdf500fb6f0b14f0c9fc43f5e901bdf016;
mem[297] = 144'hff980e85f285fd0cf9faf66f0637f9b20cae;
mem[298] = 144'h02b6f8d6ff11efaff9c7f2adf838ea81f217;
mem[299] = 144'hf37ffb74fb26fe16f2f6079d0b16f904f4c3;
mem[300] = 144'h0b43fc11f4c404ac0f81f9f7f246f4edf11f;
mem[301] = 144'hfae90441f217f4c20968fe0cf64e078fff6e;
mem[302] = 144'hed56ee160472f9ae01f0f72afb75f654fa50;
mem[303] = 144'hf6a5fa8af100f2270022ed68fc87eee8f34a;
mem[304] = 144'hf75703b10b500bd7e89200de04e1ffc4fb99;
mem[305] = 144'hf840082c08c8f0a409460e92014f0c5b0c76;
mem[306] = 144'h00e00def09690bc7f21904e4f9ed0e430a68;
mem[307] = 144'hf382ec8a06e0f8f4f09304b101c70202fd83;
mem[308] = 144'hf8820161fe820ba80271ef9af21dfc8cfd2e;
mem[309] = 144'h06b7f038faab024608def4e7f191037f096b;
mem[310] = 144'h06f6f541fb00fe6ef856080efea9092ffa35;
mem[311] = 144'hf3700e8f08ac056bf2780bc60becfed4f01c;
mem[312] = 144'h0c48f4eb037f0f8b057e0864079c008af899;
mem[313] = 144'h0947f35ff4d20b5efe480713069cefc8f6bb;
mem[314] = 144'hffd709ed0196fe17f6be01affcbffe2bf906;
mem[315] = 144'h034df5b2fdba0f6cf67dfb07ff2a0203fbd5;
mem[316] = 144'h0225fbbdf51d09810e6ffd9d0af8fc93fa98;
mem[317] = 144'h030e0ea3fb58f159f3f505b803500b29f32e;
mem[318] = 144'h00500225f1b60c80f90ee81bee0ffd65f8a4;
mem[319] = 144'hf30202ab004af2460b100b5309d205ce0568;
mem[320] = 144'hfde6f0e00694fe0ff646fe6af29d0a63f239;
mem[321] = 144'hff9804a70cf4fb380231019b08af0dc10e7e;
mem[322] = 144'hf72ff21b0ee608e3ffaa0cb8f5b4fc68088c;
mem[323] = 144'hf6e5e06ef97c001efa2ef0870280f919efb6;
mem[324] = 144'h0ca600abf194f00801f2f8e4fb31f7ccf348;
mem[325] = 144'hfaf50e11fcdb0667fa560dca0b97f06df9ea;
mem[326] = 144'hf8eb070c0b430e7ff7a5f69a0883f64bf9f0;
mem[327] = 144'hef33ff06f8eb0de20543f122f8d00327f876;
mem[328] = 144'h06d806ccf75cf2150958032ff58f004ff390;
mem[329] = 144'h067a0171ff8007320b6205e2f00a0290f922;
mem[330] = 144'h0c1ef8e3f0bff963f97004a1f836f804ddf3;
mem[331] = 144'hffeef2bbf38704aaef0ef0f7fe45037ffd27;
mem[332] = 144'h0183003a07e70353f2d9f48308b40710f52e;
mem[333] = 144'h0ee10a20f3560faff26c07550234f309f896;
mem[334] = 144'hf55ae6a8f20500fefdefeda9f536e737f0f5;
mem[335] = 144'hfacaec5f08980d90f54fed31066707c2fa3f;
mem[336] = 144'h04c806d5033cfdeffce6ea9903def6a20fb3;
mem[337] = 144'h062bff0ffb840486fb91fdfafcd4f3e2f5c3;
mem[338] = 144'h05be00e2ffa9fa29099af9caf9d3058c0dc8;
mem[339] = 144'h09b4edce09fdf3f9ee09f5b8f6c4f6d3fe9c;
mem[340] = 144'h0cb9f7b7f0c9f708f9b502f1f52bf9f00673;
mem[341] = 144'h071cfa6c05b1ffc603a40e0f04a3fcf50e5a;
mem[342] = 144'h01a90dba0e6103ef0098f63e09be0b980d40;
mem[343] = 144'hf4e404b4fecdfa0201a10b820a0bfaff0764;
mem[344] = 144'h097904c8ff03f4aaee98eeabffa10dadf3e5;
mem[345] = 144'h031ffc0200bcfb0cf9d605600ee5f62ff15d;
mem[346] = 144'h0a13e603ec7afed3fb34e7ec0199ebdefad0;
mem[347] = 144'h0677fa13026afdb90d40fb95fcb2efca0a67;
mem[348] = 144'hfa40f935f2b2f048fb90fe3e0218fc9a0922;
mem[349] = 144'h0cad0c54f812f534f56c0ad7026503de0b92;
mem[350] = 144'h0779edb5fcb7f2da09d7f123f774056a0a73;
mem[351] = 144'hf1edee51007c057d01f000d304c80b68efd0;
mem[352] = 144'hf2a8f428f2dffeebec46fedbf14306ee0bd5;
mem[353] = 144'hf97909f80d270235f572049bf2abfb25f25a;
mem[354] = 144'hf9c4fde5f5fdf91ef59ffcd30d9cf640f62e;
mem[355] = 144'hfc3ceacb0b88ef85f1f405aefe08f075f246;
mem[356] = 144'h077c044303200dbd0b900bd9000803160f12;
mem[357] = 144'hef010d9dffc60dccf17f0d89ffb2feba0919;
mem[358] = 144'h01b40213028e0b5a061008e7fb700684f7a4;
mem[359] = 144'hff0af6b0f939fbc3f7080314068ff68a0ddb;
mem[360] = 144'hf916f149006afecd03a3f313f6ad0500fc30;
mem[361] = 144'h0bc4f1820f8a03d0f5dffabdf0f1f3cb01f9;
mem[362] = 144'h04d0e4fff9c1fd6a05500a84f792ef56084c;
mem[363] = 144'h09ea0bdbfd10f1e5fa3af0df08a6055e00e1;
mem[364] = 144'hf79bfd940099fd57038c096cf5140a770bdb;
mem[365] = 144'hf7f9fcfe0d15f105f99109e6f109088dffd1;
mem[366] = 144'hfa01fb47057cef53ec2a03f7f01df05f0a33;
mem[367] = 144'h041ff3b2f17b043d03b1fc33018cf1a4f723;
mem[368] = 144'hf08effadf383fabef469fd04f9c20b68eff3;
mem[369] = 144'hffb8f255f3c90f2af1ccf6db02b706cf0f9c;
mem[370] = 144'h05a2f514014ef4d7f611f3fd03ed08a30b97;
mem[371] = 144'hfa7802a0f059efe60f010776f5340e32f7e6;
mem[372] = 144'h0a4ffd8bf9a8fe8df1e806a80088fd3bfdee;
mem[373] = 144'hf23efd55fb1e0f68f39ff91009dd0e6efecd;
mem[374] = 144'h069af267005efaa1fd480b42f9120a520898;
mem[375] = 144'hf61e0e900fef07bff1f40ddcf6da004afcd7;
mem[376] = 144'hf0d70501f4ff0dcff4f803ef0509fa3e06fc;
mem[377] = 144'h040ff918fc61f99e05adff9b08910b7f0b27;
mem[378] = 144'hf7dbf3e7f0d5fc870c17f8a8f6350bad09ce;
mem[379] = 144'h0dbf08d309b403fc0b300aa0fe73fcd0f22a;
mem[380] = 144'hf672f465fd920eef0831f2b7074d0dad0d5d;
mem[381] = 144'hf71cfbe1f47b018306d0fd2cf5c2ff960937;
mem[382] = 144'hf429feb30df4f14ef29ef6a10568f939fb35;
mem[383] = 144'hf84ffae5f01fff0a0f19091dfcb005be0450;
mem[384] = 144'h09d3f7d50231fa9e0595f6d70e9dfedc05be;
mem[385] = 144'h0401f0ddf11dfe12f4ba0615046b0400fdb1;
mem[386] = 144'h0aa000cbf7f3fc60f10ef262030cf516f82b;
mem[387] = 144'h06b0fecaf5e5ffed0145fd54f331f2150285;
mem[388] = 144'hf194073a078ffe2bf641072e0d580d4bf555;
mem[389] = 144'hf724f4cf09c70973f5730d37f14e0211fd2f;
mem[390] = 144'h0f39f1c0fa0f01690342f958fbb2f373f3f1;
mem[391] = 144'h0a190d1c014706e9037afd4e0a79fee80662;
mem[392] = 144'h0ae6ffefff74001101effcdf0866f1060236;
mem[393] = 144'hf91d0d01fa42047c0b88f7a90ec8f5d607e7;
mem[394] = 144'hee480c5dfd34ff03fa42fe240bcff94c0420;
mem[395] = 144'hf727fc2c02f4f5baefabf938fca4035efb1a;
mem[396] = 144'h0e200d7af4f8fac5041afd3d04220100f854;
mem[397] = 144'h0876013a0a27fa30020af431020dfe5ef924;
mem[398] = 144'h0891fea00e43f12c026c0712f5040476f165;
mem[399] = 144'hf67f0a2b0233f42ffff107eafdf5fdd50760;
mem[400] = 144'hf3890072fe870d56eb8bf2e1f4e2fe5c0498;
mem[401] = 144'h0745fd6d0cad0822fb12f74df3cc0a960847;
mem[402] = 144'hef6df8ccfc1ef8b3083ffef60067f150f159;
mem[403] = 144'hefadf630ffc50c790a1c0134fd930b20f3c7;
mem[404] = 144'hf2bc01010112f20c0c4407330d5ff936efa1;
mem[405] = 144'hf7dbf716f481063cf7ddff70f75bef8def5a;
mem[406] = 144'hfe8e031df9bd03e302b208df0e770129040f;
mem[407] = 144'h0320f34afe2c0ecbf0d3fbdef5130d0bfe3c;
mem[408] = 144'hf972f33b0983f61a069bf0930ca10dc70cf0;
mem[409] = 144'hf432f277f3d4fb1800d4018efbc9f25cfe5d;
mem[410] = 144'h00300d57effc06df03300416fe46030aee47;
mem[411] = 144'h05e2f6c10345f19ef71f015409b2f7b80c2d;
mem[412] = 144'h07b50361fb23fe720cf001a7089bfd440ead;
mem[413] = 144'h0f8602c604950c01f7a5f41ef4bbf7d00d7f;
mem[414] = 144'hefaff2b8f2c5f7ea0316f361fd7307bafecf;
mem[415] = 144'hfa4cfa1b0029064af65907f8fba5f3cff102;
mem[416] = 144'he2c8f60a0125fc47f247db22e3ea0db2fce0;
mem[417] = 144'h051bf4270d7b00d5eed203d60b64f6f80d80;
mem[418] = 144'h0cdc0742f5f107d2ed1701cff969f6e20d46;
mem[419] = 144'hf27cf76104eb0ccc0a59fddff643f305fb41;
mem[420] = 144'hfcff098a0447ff81f538f08d0d6c069ef75a;
mem[421] = 144'hf746f79df597f2e007780968f6190777faeb;
mem[422] = 144'h0640f4bcf12909c109a9fdadfc310aa0fa7d;
mem[423] = 144'hedcaef8fefbbfc2cf13d088a059eefcbfcc2;
mem[424] = 144'h05a9edcc02c3efd3f1f3099207f0fd6d04c9;
mem[425] = 144'hfa180200f337f26ff108f56bf8f9fea6fd8e;
mem[426] = 144'h0917fdb8f295f59c0222061b02def86f00ef;
mem[427] = 144'hf6f8ef000b720794eee8f762fb16f993fb1c;
mem[428] = 144'hf93c01e1f42ef3abf0930bca03a5f5aaf372;
mem[429] = 144'h002a0d2cf9cdf621fd5501b7079f0b640864;
mem[430] = 144'hea8be6daf0550d50f50b01befcbbf7530af5;
mem[431] = 144'hf1e3fb36fdd1eedbf2030adb045801ddf982;
mem[432] = 144'hf28e0e34f12d07da0632f143034b03f3ff39;
mem[433] = 144'hf44c09c502dcf0920ecf0ea3ff96fa300be7;
mem[434] = 144'hf403f1fa0923f8defba80ade015cfa3df205;
mem[435] = 144'h07960a1501d7faf5f3d6f5c2fb44f25f0c6c;
mem[436] = 144'h0573f85f0438fc17f41908d8ffd1f67cfdf8;
mem[437] = 144'hfa41f5ff0b040b0c05d6f892091ffaa9f168;
mem[438] = 144'h00ea0801fde3fd9bf893fa9309f50a1e0ec7;
mem[439] = 144'hff2bf64ffdea019b096b0c16fcb2f65ef2c6;
mem[440] = 144'hfe79fc96fc9104abffd3fb2afb2302c9fde4;
mem[441] = 144'hfc41feb6fb6b00faf01c01b4032d074ef8c6;
mem[442] = 144'hfc35fea0fd910698f2140c5ef9350a7dff15;
mem[443] = 144'hf5790ba606b6f6a90904f9b90bfe042efbb4;
mem[444] = 144'hf5be0f5ef84cf15a0b3ef0500a5602e2f46e;
mem[445] = 144'h029ffa130be3f94a088bf17c0016f41800fa;
mem[446] = 144'hf6a0fdf6f9f1004602bcfb5fff1104bbf304;
mem[447] = 144'hfc2ef2aefbbf0a8a0903f4aef50bf9be0c33;
mem[448] = 144'hef13f132026804ae01dff3a602990923fc0d;
mem[449] = 144'h0c2aef3af14affaaf94f064af850f6da0ecc;
mem[450] = 144'hf27902a9fe980978f3c501c2075bf481f6f4;
mem[451] = 144'hfd9aed2bffe80074ee80ee49f04405280a8d;
mem[452] = 144'hf43ceea1f907fa5307eeef8e0184f88bf0c0;
mem[453] = 144'h0450f2b5fd17f0040cd40d0ff4f9f8ef0a02;
mem[454] = 144'h0e54f9610207f11dfb10f395f106f182fbb7;
mem[455] = 144'hf1cfffbff4240b18fd60fe47f947f3fe01d1;
mem[456] = 144'hf387f150f348fbc5f09e09eb02b3063a0f3c;
mem[457] = 144'h01150e2205f00457f673f72bf2f70a520178;
mem[458] = 144'h045df49ef3d60198ed7ee9cdf6cafb41023d;
mem[459] = 144'hfccc02b80650044dff5c00b9068afeb60a17;
mem[460] = 144'h0168f34cf58b0fb8ef9a0754f04bfda8fe4e;
mem[461] = 144'h0b09f9b7f95a036a09580760f4310fe505c6;
mem[462] = 144'hf9440030ff6c09940b2ef1b1ec3f03520a08;
mem[463] = 144'h02a7f33602410b63fc7dfaab07b6f517ff9b;
mem[464] = 144'hf447f4b503ec096f000bf6460b94fc74fe57;
mem[465] = 144'hfbc0f2cc0c22fcfe0e650ee8f9caf0d6f97b;
mem[466] = 144'h043203c9fea0f619ff12f06bfd87f6ccf09c;
mem[467] = 144'h057b07c00b8cfaf0efa3ef860e4206cf00b8;
mem[468] = 144'hfb8806930042f01d06b9fae80f87f84df117;
mem[469] = 144'hf8c40d140db7044e0661ff7e0a44ffb0f1bf;
mem[470] = 144'hf3a4fe38fac409540b59f81dfd3700f702a6;
mem[471] = 144'hf3eafdb1f041f39ef0f8f8a7f35208f6ef4e;
mem[472] = 144'h07b10186fc89f6ebf374f9c2f138efe1f759;
mem[473] = 144'h03820f15f670fbd2f6a3f122f596fb41093c;
mem[474] = 144'hf74008c9f3ef00950ae602dafad5f56507d5;
mem[475] = 144'h066a0cc6f7250897fb3bf628073d00ff08d3;
mem[476] = 144'hfe2a0b9efcd7026ef162043708c8f2750401;
mem[477] = 144'h0095036ef822f50d0081ffc3f681008ef454;
mem[478] = 144'hf699069df81b093ff41d03a2f8b702050aee;
mem[479] = 144'hfe840c1af08ff424f0c40e1b07c50323f9cf;
mem[480] = 144'h0e1d0367ff3bf8b808d406d20c18f9f4f0a8;
mem[481] = 144'h009efd6d0b10f707f0ea0837050805b406ac;
mem[482] = 144'hfa4af29306fbfb5affdb0772f2800faef417;
mem[483] = 144'hf45a07900531ffef0ef7f30ffd240be5fe64;
mem[484] = 144'h0cd809ab0961087cfedc052301da0609f147;
mem[485] = 144'h0c18fd7a08fcfe1bf13cff350f950209f577;
mem[486] = 144'h0e2dfe56ffdf0914f69b04b1f0660f49fd88;
mem[487] = 144'hf498f877f5cbf275054cfab8f7abf91c0c5e;
mem[488] = 144'hf9c1f224f69cf15d04ec0608f2af0a12f715;
mem[489] = 144'h05880a47f43b0310f85ff27efe5202080042;
mem[490] = 144'h0513039a0ace075c040001f8ff8608e1f62e;
mem[491] = 144'h0b8f07f0f47a0822f154052f006c06c0faea;
mem[492] = 144'hfc6b0ce10859fd5bf663082b0a7ffb4ffb73;
mem[493] = 144'hf1180870033001e300e4fab70d9005e00b1e;
mem[494] = 144'h054cff4e0bba04b00d94fec9fad1f3f0090f;
mem[495] = 144'h094904bc0019f32c0d0ffa49054ff0c00051;
mem[496] = 144'hf925f952f522f90005eafe29f1b2fc1efd9a;
mem[497] = 144'h0fa0f7850233f75efcb400ccfffff9270cd5;
mem[498] = 144'h0f420b11f418fb0c0b8ff4d20dd8038f05c2;
mem[499] = 144'hf5cff938fa97f2d3fb4d0acd087b0349f4c7;
mem[500] = 144'h0eb9fc0205b20f0ffb6d02a2039cf55604f8;
mem[501] = 144'h03840fe60a7ef0690e32f89c01f404810fa3;
mem[502] = 144'hf43bfab1fd2105baf464f284fc34093ef0f0;
mem[503] = 144'hfb480d00fcab0af4f1abffc209e801d0f1cc;
mem[504] = 144'hf37a0622fa25fee3ff7604a305f80411fd65;
mem[505] = 144'hfc94fff107dffdfdf3880abafa64f8000fda;
mem[506] = 144'hf3ddf2bbf6db07c207bbf92fff59f02e0ad7;
mem[507] = 144'hf270063cf0180d27004b0356ffa4fb3408d7;
mem[508] = 144'h0065f941063509960a7d0700fb73f8550de8;
mem[509] = 144'h0ccaf6f303e7faacf9c7f5bbf1810266fb55;
mem[510] = 144'hf43d02c802b9f4cf012b0076047d07910971;
mem[511] = 144'h0915f24afb32f0d0f3110095fdbf0b12f5d1;
mem[512] = 144'hfef7f363081106e0fa030a50064d0681f35a;
mem[513] = 144'h0e700e8dfeb5fdf8f8bffdf2fe13f0eb0bf7;
mem[514] = 144'h04d40b7e0e6702ad020bf263f125ff48f0e4;
mem[515] = 144'h064d037ef9f3f894fde0f296062ffdd7ff38;
mem[516] = 144'h07bef9970e9ffb7df3f508c9f480006ef086;
mem[517] = 144'hf548fca9f8c4f4a40de0033cfaf40168faea;
mem[518] = 144'hf3b10616f8e40e610b9a09c4fd12f776f88b;
mem[519] = 144'hfd54fa1af4d0fa400952f432f7db0bdef5d1;
mem[520] = 144'h0eaaf32e0a7b020cff9a01560cb40f90f60e;
mem[521] = 144'h0cd60ac00d8ff5d0f778fbe1fed40bea059f;
mem[522] = 144'hfde30065fceef63efa20f7bbec14023bf147;
mem[523] = 144'h0139f1e0025c0ca80c8e08c5f388052cf153;
mem[524] = 144'h036c01f1f6c7fb7dfbc005a0f4cafc580649;
mem[525] = 144'h01aafe6c09eff4a707a00488fbcff9f707ae;
mem[526] = 144'hfb19ff7ff92ffd0d02c301720aeb03f9fcd6;
mem[527] = 144'h0c960b8bf46df6e00498f30cfac802db04f4;
mem[528] = 144'hfaf8ef2b092ff2e0f6d8eaf90428f57cf111;
mem[529] = 144'h0935fae5f1b30ce5fa4a032af997f8d50a7d;
mem[530] = 144'h0ab906de06fdfda4f418efe2030bf61d0a29;
mem[531] = 144'hef3d00d1050bfab5f72aef38022af5ab00f0;
mem[532] = 144'hef170982036ffca1f058efb5f79ef4e80a61;
mem[533] = 144'h0cccff13fb1202c3f02f0bea0e38ef4e0009;
mem[534] = 144'h0c33032c0a2dfc85084401b6012efb9ffa68;
mem[535] = 144'h08d6ffcf03cafe1b02d5f002f42b0a03f512;
mem[536] = 144'hf84fefa7ff6d05c5f79309e2f8b9f022f413;
mem[537] = 144'h00880b480ebcfb5cfc22fe7ef05deffbfc7b;
mem[538] = 144'hfbd1084cf9f804e2fd03fe7afcfaf105f90c;
mem[539] = 144'hf8c9063f000702370102efc10d6a0df50182;
mem[540] = 144'hfca3f7fef08001f4fd60fe09f020ff7a059a;
mem[541] = 144'hf08b0b2ef26e05d8f81f0282f0b5fdd2f761;
mem[542] = 144'he045f70fefce04dcfc28f463ec05fee300a3;
mem[543] = 144'hf4fe0576014209d8f23902e8084efdbef085;
mem[544] = 144'hf4d50cfdf89e0a39045b0977fdeafee40139;
mem[545] = 144'hfbfcfe93fbebf9170885f97d01c0f38ff119;
mem[546] = 144'hf3090cc602c7ef040a78f0b305a30cf7f78e;
mem[547] = 144'hfb9608b0f4ae084bf4c905af06f8fb85f9e0;
mem[548] = 144'hf9a8fc17f64d0af9fedef20606c6f3c7f4ec;
mem[549] = 144'h0095f1e50c100b98f232fcf802c7fbdc0d2d;
mem[550] = 144'h0d81f2cdf08ef3b0071b06720ac7f28c09d0;
mem[551] = 144'h0be1f040f2e004e2fa9709890c6ef9f3eefd;
mem[552] = 144'h0d3d0ae9f30e0dd8f2d9012cf330f94bf7d5;
mem[553] = 144'h022bff0a006f0d5007c50aeaef5600da0085;
mem[554] = 144'hfa3307fb04f6f398f8d7f0d1fd1bfcbe0a39;
mem[555] = 144'h0853f09af96ffd00edacf2700b33f808f31c;
mem[556] = 144'hf7490bf7fc090e38f0b606c4f276084a0a44;
mem[557] = 144'h0dcf0391f343f70b0b6a0fa6017af0cbf4c8;
mem[558] = 144'h03110208f775fdee0a3a0913019e01830c6d;
mem[559] = 144'hff5103dc0ce8f89cfe550862015d081af81b;
mem[560] = 144'hfaedf5c4ffc0f368faef02feed37f27f0322;
mem[561] = 144'h0628f7410739f84afda6fd54ef57f2250cf5;
mem[562] = 144'hf22a03f80157fa6102cff4cdf1150546fcf7;
mem[563] = 144'hf3b8f01dedf1f34afa07f642fc56fb11fc1d;
mem[564] = 144'hf2fe0a6afca2f2830d20ff8c014d05bff601;
mem[565] = 144'hf21dfc7cfd820364fab20b50fd1cf632f0dc;
mem[566] = 144'h04fef16c072504c002720430fe0ff21dfbbe;
mem[567] = 144'h07b1fd110adefd5df285f0a10232eef8f3c7;
mem[568] = 144'hf26cfe13f3e8feff03b8f8d8ed860dc5f8c9;
mem[569] = 144'h0f93fff903eaf47000c60e65f063f4f3f6fd;
mem[570] = 144'h050700680658f2adfe12e7cdeefcf2c0f372;
mem[571] = 144'hfa53f6cf0d620a55eff50289001cefcc0d6d;
mem[572] = 144'hf82fefea0b2d023cf98e0796f918fb79f820;
mem[573] = 144'h05c9ff2e0df206b809fe060f0c6d0922f1f9;
mem[574] = 144'hf6e4f9f00ac2f5bff8cbd90af6b9f59efd87;
mem[575] = 144'hf763f3cff60e0a6eecf6ed3af68204ce0943;
mem[576] = 144'hfa63f700f71d0e18ec4afc9cf2a4f4120763;
mem[577] = 144'hfd3e024a0084fb48f1750507016502900414;
mem[578] = 144'h0e020fc6f72c00bfff31fbb0088805e104cb;
mem[579] = 144'hf8f9f0fc012dfbf90466fd5df56b01eef567;
mem[580] = 144'hf71004c1f7720e43f6dff562f4890ce4f2ab;
mem[581] = 144'hf9a00d9cf83d0ccbf38405d50702058cf57c;
mem[582] = 144'h01a8fd7d0e5d0c45f9a40e8507b7fa080dbf;
mem[583] = 144'hf06a04ef081ff92a02d1f4cff0ab09dffbfc;
mem[584] = 144'hf84ff0080800fb2def12ff10f13308a4fcf8;
mem[585] = 144'h0f3bf45a01a70f78fe70093606b40a9bfa4f;
mem[586] = 144'heb8302f1f228fee9f83908bcf8ccef05ee95;
mem[587] = 144'hf063f0d103760d17f8a2018c0cd1fcbef65d;
mem[588] = 144'h0c1a0a96f215f214f26ff68a0eab0e96f621;
mem[589] = 144'h0371f93a0488fc4b01ec078c0d3af8d207c0;
mem[590] = 144'hf918fe3dfa05f0cdf1ab029fec97fc42f467;
mem[591] = 144'h0152009400570430f58c03c4fb360f0b0170;
mem[592] = 144'hf94a04a4f5c006b90a47f4b2f6060df5f7e0;
mem[593] = 144'hfbd3007dffc8ff88f15509e70da8f03a024d;
mem[594] = 144'h070f073e0c36f1930997f8760cfcf56a0d61;
mem[595] = 144'hf30afa1e040e0d28fd32f7560baa07020a59;
mem[596] = 144'hfca1f387081e004ff270f2830138f6c30d18;
mem[597] = 144'hfa6ef01607130706ff33feb5f7610414f500;
mem[598] = 144'hf49f0d42f9f4f4ed03dd0ed20507076200e8;
mem[599] = 144'h0cecf13afe37f01d09c70488fe82f6ecf53c;
mem[600] = 144'h0e12036703d5078cf4900b760c6706a0f634;
mem[601] = 144'h018104350c2ef617f4320049092f085b0a61;
mem[602] = 144'h00c6f0a8fa4100650893f6c4f920ef8b0286;
mem[603] = 144'h0e2bf98c05af0ca40c52facf06e5fa26fc6c;
mem[604] = 144'hf3c1f043f28bf4f0fda8032d0b25fac9f385;
mem[605] = 144'hf6a3f5d3008ef99306350cc4f47efbeb0ded;
mem[606] = 144'hf8cbf6e505a20e64f4ea09aef8a60796f86c;
mem[607] = 144'h0944f5eb08600117f43cfd200812f17cfb29;
mem[608] = 144'h04e1ef8b09d9f44bf37900e008e7040c073d;
mem[609] = 144'h06a10f4b0a900a0800fcfa35ff690afb079f;
mem[610] = 144'hf0b7f1d10071f6d2f930f4c20209ff07f953;
mem[611] = 144'hf1b6f6b50721f7f4fd3202220ad60fb50578;
mem[612] = 144'hf74ffe870090fa7c0035f6c203f2f565f524;
mem[613] = 144'h0241effa01bffc1d06dffc6a09f8fd6208da;
mem[614] = 144'h064af36a0bb3010407f4067009e0fd3106f5;
mem[615] = 144'h024e0233fd6ef02df382f9e6f238f1caf11e;
mem[616] = 144'h0c8ef7d80658fdaaf53bfea3fd840762fadb;
mem[617] = 144'h086ef670f0a7fc98f98d0af8f65ffc4208a8;
mem[618] = 144'hf066f0380ebd06eafb1b0a76ef1dfe6b041e;
mem[619] = 144'h0d1009fbfeddfc84f5fa0879fd89ff5801e9;
mem[620] = 144'h088e0002fd9f08730dac08ddf193fb2e0036;
mem[621] = 144'hf258f4f9077df7350eeff9460428f8c8fd33;
mem[622] = 144'hfc84fa5b0e11074afb62efd0fa200951f223;
mem[623] = 144'h0d89f18ff4370d12f239f8ef0559f18ef64a;
mem[624] = 144'hfb8cf220f1d40b170a7efe52fc7bfda6067f;
mem[625] = 144'hf72204edf054f71807d8046bfa02f1fd0031;
mem[626] = 144'hf300f01dfd4608200b5a037bfd9509710ec3;
mem[627] = 144'hf227effc0d9806d0f6e9fe70f03c09c5f548;
mem[628] = 144'hf4dcfa28f32fff57f95501580563092ffb0c;
mem[629] = 144'h05430051ffebfb150336fb9efe030bacf0ad;
mem[630] = 144'hfc8cefdef9d2fead0bdff35e0f3f0ad1fd06;
mem[631] = 144'h0ba5fd920ca1f195070d0a80fb950a0ff489;
mem[632] = 144'h0494fb860e6d03460ce3fd71fccef2a6ffa0;
mem[633] = 144'hf7990d7efae2fc72f1a303a50cdd01730d7d;
mem[634] = 144'h06c8fffaf4fbfa8dfeb4fc3cffe40d32ef37;
mem[635] = 144'h0d1f08130f420a56fb9c01c1efbe0a47fc6e;
mem[636] = 144'h02baf48ef528f16907c0fef9fb4608e8effb;
mem[637] = 144'h0da302f2085dfbbdf50005f70c3f0ac10f38;
mem[638] = 144'hfb1608f0f8bc0988fa8b08340e130ecef649;
mem[639] = 144'hf41ef9040e19ff5d08c4010dffca091c0568;
mem[640] = 144'hf39cf997f6170dc5fab4fbfe0a530669000b;
mem[641] = 144'hf57f0af3f868f0a403800000099eff790baa;
mem[642] = 144'hf3640a8b08ad041900a0f33b090ef34408d6;
mem[643] = 144'hfc04f41ef919f99a0b48070ff196f8d90369;
mem[644] = 144'hfd8209b205ad06840896f2a205820384f268;
mem[645] = 144'hfe0108aafaed0d87f2fff4cd07200210ffa6;
mem[646] = 144'h0272059af79af8d4fc1e09da0a3b029cff9f;
mem[647] = 144'h0bd7f00bf953f162f68d06aa035df28bf267;
mem[648] = 144'h0451f8fdfd0b0a83067202bf010e0be10d4a;
mem[649] = 144'hff7e0f6af452f1da091501650c77f2990c9a;
mem[650] = 144'h07ea0595fb53fe76f81401d204ed06f301df;
mem[651] = 144'h089106cdfea3fcb8fe9bf668fa86f553f85a;
mem[652] = 144'hfaf6fa2503bd07e3ff090e23f5ccf253f75b;
mem[653] = 144'h0883f0eaffa7fe8a055708c1f9e2f199facf;
mem[654] = 144'h0d52f7a30006ff0f0b38f7c40082fce8006b;
mem[655] = 144'hf3a9fccb09eb0e96fc590247030d08e3f956;
mem[656] = 144'h0733f6b80f2800c6f6b0e975f039007c0c54;
mem[657] = 144'hf6e9f1f6f446f8f70c8ef3faf43df510f477;
mem[658] = 144'hf751f9b1060e08faf0fe05bcf79a08b0f293;
mem[659] = 144'hf7a9f447055dfe280a1eeea002bb089a05e7;
mem[660] = 144'hf586febb04d6f55ceebef0f9f7e607c702e6;
mem[661] = 144'hf83ff75fef60fc34f9d5faea00def75e071a;
mem[662] = 144'h0ec306fdf71709b3f2b10672f5eb053e0193;
mem[663] = 144'h06d707d6fe23ff5804cef0620b43f47f08ec;
mem[664] = 144'hfa66f3d6f698f24bf226efd908310ad50d54;
mem[665] = 144'hf0c50cbffd46f7edf9d2fedb013b01dc0c84;
mem[666] = 144'h07eeeae2f3d408b7ede7f4110608fa87f263;
mem[667] = 144'h07d403f10ee5f03a04f60e61f4cbf77a07aa;
mem[668] = 144'hfc78fb7ff544f16ef6cb012207dcf74ef071;
mem[669] = 144'hf525ffc5f06e08f80502fdb6fce40259fb84;
mem[670] = 144'hf41bffc0f65908f4014b078bea8afb6a0625;
mem[671] = 144'hffb6fb650cd1fcebf112fcf6f834074afc48;
mem[672] = 144'hffaf05f90237fcae08d4f7b80725049e08cb;
mem[673] = 144'hf8d6fd76f0f0f96a08bdf9aaf260fd7604fa;
mem[674] = 144'h0b46f8800fadf06cfec70ba30ed70b57f599;
mem[675] = 144'hf5230d37f76b04dbf9460e16f74f001ff094;
mem[676] = 144'h0d05f2430c7c01c2f7b40dbdf3f10145fc1b;
mem[677] = 144'h07220c9bf8e7f045f26ef73401a3fd9c086d;
mem[678] = 144'hf04bf789fb5afd8c079f0d850baf00d300fa;
mem[679] = 144'hf4d801200ad0f78403e9068207e7f11ef55b;
mem[680] = 144'h0581f3a9f4fcffdff933f05dff59f1adfd8f;
mem[681] = 144'hf3f6fff2045f0023fecffcab054dfbc50b46;
mem[682] = 144'h04b2f74ff80cfbf20972f142fade0875f1d6;
mem[683] = 144'hfba80bfb0dc7fd09f743f99bfa6cefd1f656;
mem[684] = 144'h033e0a040766f60cfdaef0f3f059f93ef7c7;
mem[685] = 144'hf55ef1b00a1af0f5f83d031af3c0fe14f205;
mem[686] = 144'hf3e0fd6af7fcf30704430721f8aa03a80776;
mem[687] = 144'h061a0ad2011cf9a70ac404a5f853f84ef657;
mem[688] = 144'h0017065802a9fe21f487fabff4cb08e5ffd4;
mem[689] = 144'hf14cf153f9420a6e0828f35cfe400b9e02f9;
mem[690] = 144'hf383f37602f7f05ffa4cfe250f84f317f616;
mem[691] = 144'h03b5047e0cbb05de0f07fd42f0a4f03a00aa;
mem[692] = 144'hfc0bfe8affa803c4054900420ed3f965ff13;
mem[693] = 144'h0f7b02810b0cf2cf0a0809ed0c68fcd0f9ce;
mem[694] = 144'h03e30c35f5e5f23af576f31df43bf2f30003;
mem[695] = 144'hfeaff09af5d4fb97f6610633028c01fd0b21;
mem[696] = 144'h00a0f223f4610a130615f963fcb808cefd1b;
mem[697] = 144'h0af4faeff00ef2bf06320fe30ab3f1c60f50;
mem[698] = 144'h0548068cf28b0624ffaf0318f78a0ec6f399;
mem[699] = 144'hf733f429f46102550ab903d305f804bb03aa;
mem[700] = 144'hfdde0a7e0f6e0d5c036606e209ae0fa703ef;
mem[701] = 144'hfe4bf6390ee30a9e010505a6f213ff0c0bea;
mem[702] = 144'hfa1bf1b80396fd56008f052ffae90b530c47;
mem[703] = 144'h014f0e58fefef315f3ccff1809bc0312f903;
mem[704] = 144'hfa520b410e63066e032ffbd90ad003c2085e;
mem[705] = 144'h01a403430c9af454fa590bdcfee50501006d;
mem[706] = 144'h025cf5d0f500fcb2011bfcdf00f8f21af32c;
mem[707] = 144'h032cf3580555fde30bd5087302570822f82c;
mem[708] = 144'hfb4c0e9efed3f4daf63e0f70022102d30f93;
mem[709] = 144'hfe360adafa0b068c0fa9f9c8f6d1ffccf647;
mem[710] = 144'hf47b02fd020ef4a9087b085bfc4cfc82f175;
mem[711] = 144'h03a2facbfc200b7500fe0c6605640c01f788;
mem[712] = 144'hf7e3099ff410fc1ffe3407c1faf8f3340fd8;
mem[713] = 144'h0b6f0ab100400a46f5bc08e307ddfd1eff1e;
mem[714] = 144'h062b00a9f2a3f68b00a4062bf4a8f35508e3;
mem[715] = 144'hf3d4fc2ffa4bf60bfc920713fa8405a10e19;
mem[716] = 144'hf0b3f626f069f097fd9f06160db0fe920b5d;
mem[717] = 144'hfbcb02a4f650084407e00c590747f442034b;
mem[718] = 144'h02dc014a0336f2b00a840bbe046ef12e001e;
mem[719] = 144'h0598ff49f2d7095b0d090ae3fce9f36d0a8e;
mem[720] = 144'hf63901cff32df8520dc2f490016afff00550;
mem[721] = 144'h0e23075ef5360a0f00b005b5078f0eccf7d3;
mem[722] = 144'h0d74fc44f42ff6a30e5bfd020c80f1e00d1d;
mem[723] = 144'h02aa096ef925f0b30a1bfd73f0db0b0b003d;
mem[724] = 144'h0f5afe3a05300e720fbc06f6f68af538f538;
mem[725] = 144'hf65bf0020e1f0cb7044301ce0362fce3000b;
mem[726] = 144'h098a02c20afc00c405b5fc29f43afe3e0af1;
mem[727] = 144'hfea4038ff2310d7cfe8f0d1f0f62f95ef819;
mem[728] = 144'hfb06fe66034ff441f09908450c6f089a0ec6;
mem[729] = 144'h0f7cf28ffc51fec7f34a0682025300080e0a;
mem[730] = 144'h09b1f449f48ff0b700e4fce30a44f940091e;
mem[731] = 144'hf963066c08b5080202420422f565f9f0fd16;
mem[732] = 144'h0167f0d8066d07f3f81b0c300aac049201b2;
mem[733] = 144'hfa5ffa50057ff5780baffb96059af782022c;
mem[734] = 144'h02780867f3ea08a4f435f85dfb18f369fd40;
mem[735] = 144'hf302ff21ffbd0af20126f9f608a605990a60;
mem[736] = 144'h0b1001ff0bd7f0e9044dfa100e5fff490f25;
mem[737] = 144'h090405b80f910b8e04820a420637fca40f24;
mem[738] = 144'h0f3b0ac0f56102cdfba70bcbf75dfe74f188;
mem[739] = 144'hefd70665f9e8fcfe048709b7f2c9f6b80f0a;
mem[740] = 144'hfa15f4d10dc8f6870801067df840fbb10e05;
mem[741] = 144'h047a0466053b0a8df990f8eff6770b3cf0e5;
mem[742] = 144'hf247fd05fe47f924f6ecff780eccf19f09c0;
mem[743] = 144'hff55f4300ba10e2d037df9bdf45a04620ac3;
mem[744] = 144'hf54602cd0eb4070bfaa2f28cf84908c90a12;
mem[745] = 144'hfad2f2abfe0f04af06cbf99dfc84f33f0fbc;
mem[746] = 144'hff0800f9f09cf04d0a96fb99034e0790f114;
mem[747] = 144'h07d9fbcfefd9fd19f4b0049001860d36f095;
mem[748] = 144'h0972f116f1fd0f3d0053f60ef2c90e6efe2b;
mem[749] = 144'h0b96f084f63ffd1a0accf903ff13f4dff8cc;
mem[750] = 144'hf4420e4505bcf848fdca08370f5e05df0722;
mem[751] = 144'h0033fe61f4d30374f090fe6dfd34064dfdce;
mem[752] = 144'hf87b00e40c800e50f187f8fff268f379f3bf;
mem[753] = 144'hf7b9f1f3f43301b1005c0e46010ffd2e0d51;
mem[754] = 144'h0cf0085ff21b0a53f0d800ddff4e0c230d1d;
mem[755] = 144'hf7f206d906eb0ae40ab8ff82fb8bfe620a2d;
mem[756] = 144'h0c8c02a8fa740c0bfa82f967f2e70cddfec8;
mem[757] = 144'hf525f84df053ff850b5409ca08780d13fdb9;
mem[758] = 144'hfa8ef2810081fe68011e01f9f27506f1f1af;
mem[759] = 144'h0603f075f304f05ef610feedfa5af725f7d9;
mem[760] = 144'h05fdfaabf5aaf3280911f9c4069cf10f0513;
mem[761] = 144'hfbcc03e5f406f67af4f1f911f15df51af55a;
mem[762] = 144'hf705fb220ba00f7cffbbf65df06b020cf0de;
mem[763] = 144'hf1b906cb0e03ff99fd7e02dc0880fd1f0021;
mem[764] = 144'h01cafa33fdd5f29e0b4c0cf7081a0523f826;
mem[765] = 144'h0144f7060db10d50018ffbd00f68fce5086a;
mem[766] = 144'hf051f893002b03fdf445f28efbed08010900;
mem[767] = 144'h04780993ff79f2cff250f9e409b90c56f3f3;
mem[768] = 144'h010c0b21f6c60fba06460a2c0dcb0d500bc7;
mem[769] = 144'h063e059dfef4f064052b042cf69a08ee04dd;
mem[770] = 144'hf10d0f49fbf2076006f9f3780c83fac8f3d9;
mem[771] = 144'h04bdffebf4c00d0ef0eb00e1eff70c230b54;
mem[772] = 144'hfb7c0e28f075f755013e0e3605acfd150e13;
mem[773] = 144'h05ac069b0758f8280d36f55e06c80516026c;
mem[774] = 144'hf7dd06e706dc09520354f340089df96e0c83;
mem[775] = 144'hefeb0180ffff0d3207eaf388f327f084f648;
mem[776] = 144'hf552f61df19f07f0fcfdf666fe97fcc0f06b;
mem[777] = 144'hf998f402f7930c10005b0224f17b0ac20d4e;
mem[778] = 144'heb2f0822f7b7fac603faf3e6f9b1ff71f46a;
mem[779] = 144'hf2fdf3a1fe2d0394017ef9bf007ef7cbf058;
mem[780] = 144'hfc42fba60b8c0adf0c32f21eff2405ec0f90;
mem[781] = 144'hf25b02b90d6305a50e32000df8750b240373;
mem[782] = 144'hf617f199fa3df48af234f934fafef653f9d1;
mem[783] = 144'hf410fa940c0af832f355033cf2bfff010e4f;
mem[784] = 144'h014cfe1ef53208c1f805fadffb55fdbc0204;
mem[785] = 144'hf04af9cffbc5002ff75f0063f4df0cd2f384;
mem[786] = 144'hfcd806b0073e0d87fa06f66304d4fdd7fb4d;
mem[787] = 144'h06a3fb6ffd910261026ef009fe99f2980c82;
mem[788] = 144'hefa60aa208a8fe8eff30fce20df50a63fa7f;
mem[789] = 144'h01dcfa63fc19fea3f1a6f05c054afbd8f226;
mem[790] = 144'hf21d0b0b06ef0a610b7bf2c108920f9707f7;
mem[791] = 144'hf217033f0090f8aef99ff273f280040b0878;
mem[792] = 144'h0b6f0181063306470781f0400339f5ebfc34;
mem[793] = 144'h0fa20f3fffce0a9200b1f442f98f08e8fc1e;
mem[794] = 144'hf958f2ae046a02f3093ef4670ae50731fea5;
mem[795] = 144'hf6830e29fead09aaffcbf130f1840248f802;
mem[796] = 144'h068a09710dbf0ed005a5f25cf917fea1ff8a;
mem[797] = 144'hffd1018ff980f1080fe903830375f21800a1;
mem[798] = 144'hff5e029c0821f803fc5f007105aafd140c30;
mem[799] = 144'h044a0723f06ef6880479082dfb900bf50eba;
mem[800] = 144'h0635f95c049d0df8fc9f04d0f07afd5bf3be;
mem[801] = 144'h082afa6604cd065f0def0178fc9d05660074;
mem[802] = 144'hf75af94ffbd000470419f3c5fc8ef328f69c;
mem[803] = 144'h0232f4caf6db0a4c0bd9fc81ef2bfd95f8c8;
mem[804] = 144'h067df081f1bc0ccdf65af1e0f3a50e700bdd;
mem[805] = 144'hf83ff4150ec5062205c6fae3fe300aea053d;
mem[806] = 144'hf7aafa7bf14f0275f0a4009cf996f2500cfe;
mem[807] = 144'hed4201e9ff9df29df1c8006d01aa001cf811;
mem[808] = 144'hfaae0a5af2260ba3fb9b028a0b2e022bfc7c;
mem[809] = 144'hf3fff252f83af35dfcff07510687fbe60cb5;
mem[810] = 144'h01cff357f497f9eb035904bdf72bece6f89a;
mem[811] = 144'hef640dbbfc56f4e30a480ac20dd6f531f48e;
mem[812] = 144'h00650bac08d8f71a04fefc44fd500421077c;
mem[813] = 144'hfa1f08df0086f22f068e06d6f79cfec5f300;
mem[814] = 144'hf695f403f05101c4f043035af4eff851091a;
mem[815] = 144'hf2700b6df307f905fef305e5f65e0598f7f6;
mem[816] = 144'hf73b0293f568ff7ffafcf7cb0e89f0ba0ecb;
mem[817] = 144'hf9f607150bdd061af28a0f78fdbbf567ff62;
mem[818] = 144'hfcea00c5f0d1009ffee9fa870a59041601ba;
mem[819] = 144'hfd94ef78f4fbfaeaf6a4f4fb04d9f6780be7;
mem[820] = 144'hfc340a92005e027e090df114050f0162f0c5;
mem[821] = 144'hef87f9fef60007de08bbf33af726f4c50b97;
mem[822] = 144'h00120b9afc9508e501c3f292fcb1f00cf125;
mem[823] = 144'h093cf93bfed2098e0229f2d1fd990e580845;
mem[824] = 144'h05aefd6bf7f50aa304a604de03c7048ff288;
mem[825] = 144'h0f4f01cbfec8f53ff3a8efd8f9330973f0e6;
mem[826] = 144'hf8fc09cc09cafcd4081506b4066df5880734;
mem[827] = 144'hfcb102b1ef850f7107a70480f0c7095009fd;
mem[828] = 144'h036508a10837f1e00e70063bfd80f1b20062;
mem[829] = 144'hf6870ca2f432014e00e9f07501d0f0eaf8a6;
mem[830] = 144'hf77f0b8a0851f022f924fbfbf33df451fcb7;
mem[831] = 144'hf0dc08fc0722f864f74605340975f60d04f7;
mem[832] = 144'hf543f96cf3a5f3d000f907b2024f001c0aba;
mem[833] = 144'hfa30f35ff95a0c5afcef03f20f1cfa34f22b;
mem[834] = 144'h0d0b07acf02804ed0ae4fb52fc5400e8023d;
mem[835] = 144'hf3cff434003f0ac8f28c04ea0391f20bf7e9;
mem[836] = 144'hf3970d3a092af0fc0414fc6508be05380692;
mem[837] = 144'hf6c6efdff4a10f45f1c6efeff5cdf2f5f162;
mem[838] = 144'hfc6c0a1b0c71fb45f2b8f46b0167f6180037;
mem[839] = 144'h02f109ab017103faf785fa0e0be9fcb70c36;
mem[840] = 144'h0a5f09fef02afa100c3f081f045cffbe0fc0;
mem[841] = 144'hf385046df693f6f3012cf060fb0209a807d2;
mem[842] = 144'hfeb5fed4fb9c098b0543f2c606ad0836fac3;
mem[843] = 144'h0095f9e7f647fc300cb10dc4feae051dfd49;
mem[844] = 144'hf20802fbfa620039fe99f2a8ff0f0c1af20b;
mem[845] = 144'h05c1ff5df36603b708e2fee9f984f2e3f27f;
mem[846] = 144'hfa990ba80df9f13e067bf4e60aaefb320875;
mem[847] = 144'h08b30cb401defd94f2d60b9c025003f9f84e;
mem[848] = 144'hf8d6f306fb65fe7af69102d3fcc00e8af1d4;
mem[849] = 144'h0831f7f0f8a105ee0edd0b070d6ef8a6fc6d;
mem[850] = 144'hf9070d9904dd0b23071e0174fedc072af98c;
mem[851] = 144'h0718f18409d40be0f6f4ff7600d9fd6cf576;
mem[852] = 144'h0ab10f440137f878080402c40c9d01110b19;
mem[853] = 144'h044fefa5095a069bfdcffc400137f436f21a;
mem[854] = 144'hefebf5e6018cf0dbfa850bd7fd9209970305;
mem[855] = 144'hfd06fc07f5e8019b05a2f9d9f4480df6f5d6;
mem[856] = 144'h0b150308f238f29607bf0a590de5f7b2fc6c;
mem[857] = 144'hf630ff16041e0f2af28af9fa0167070bf585;
mem[858] = 144'hf0dcfb38fc95f9fc0d550a1ffb4a0ca3fa22;
mem[859] = 144'hf6bff886025000e9ff39f2ce0799fbd4f600;
mem[860] = 144'hf47709350de10ede09f5f2de0298fc74f815;
mem[861] = 144'h04c20e9e021bfc9ef028f0b2f3f3f398f113;
mem[862] = 144'hf717f0b9f5750d78f8eb03870aef0340fcf0;
mem[863] = 144'hf90f08c901370daafe6aeef40d78f7b100a5;
mem[864] = 144'hfc86faa0fc86074a0a13ea41004df837f866;
mem[865] = 144'hfb28fd41f1d70d56ff16fea1f8b7f733099f;
mem[866] = 144'hffeaf30b07a3f46afaeaf2dafc9bf2ff0804;
mem[867] = 144'hfbc1ff52f76f0357f8b5f396fe09edd5f4c1;
mem[868] = 144'hfc4a07910855f7970739ef7bfeb90653f85d;
mem[869] = 144'hf607faeb0e13fd2904c70a5c074af8f5fb0e;
mem[870] = 144'hf34d0442fc360b1a07b5f7c4f31bfe0af09a;
mem[871] = 144'h0c050a6bfbb7eedf0c57fe98f1010dbb08ca;
mem[872] = 144'h0d5e04cffb1c05affdac03b00d58f604fd65;
mem[873] = 144'h04a50a9c03d507460ded0abaf514fff9f525;
mem[874] = 144'h0e3f0d7af4a1f0def420ef94f486ef21fbd8;
mem[875] = 144'hfd38030a00ab0196fe76f427f57efcc408a7;
mem[876] = 144'hfffffe23f546faaaffac0a6201ba0e6702d4;
mem[877] = 144'heff507ac043cfec8f28ff833fb5afa5cf717;
mem[878] = 144'hf9d5e921e8df0669f572f8c201fe070df318;
mem[879] = 144'hf1b0f9ae09f6fb450b26f9180145036cf387;
mem[880] = 144'hfb0af694f284057cfba905f9faa8076afce1;
mem[881] = 144'hf678028ff5e5f015035ff04b0b7006590926;
mem[882] = 144'h09b4f6e9f1db05d7ff620582f99a0c01f05d;
mem[883] = 144'h0b0cefbd0351fc4400c2098efdaaf6e10b2f;
mem[884] = 144'hef4af7b0f962f690f3b3f957fbf904310387;
mem[885] = 144'hfd750b220d11ffdbf1fcf51201630998f5b1;
mem[886] = 144'h0d02f2600f46fab701850af307ebf983f2e7;
mem[887] = 144'heff3ef09f5b2f930063b0469f95ef5370b86;
mem[888] = 144'h0a83f30b0bf2f24cfd72050a042df7900ca0;
mem[889] = 144'hf85efbb20f4ef8840c65fcd40242f043f463;
mem[890] = 144'h09d105fdfabaf539fcffef110885f0b0f418;
mem[891] = 144'h00380c8afbbbfc97faf8fad2fcf6f02f03bd;
mem[892] = 144'h08490028f141fa760ee5fc2cfaa50476f074;
mem[893] = 144'h0c160524f4f5fe8d060e046c0291f75c0ed7;
mem[894] = 144'hf8900be4fa39fd1ff02efd7302080460ff35;
mem[895] = 144'h0babf9750a58f170f19d0c78f2810db6059d;
mem[896] = 144'hf712045205ca0bf6f27ff056f6cbf3a303ff;
mem[897] = 144'h01fcf9c6084e0a33f04bf79601e4f9e2f3d4;
mem[898] = 144'h0638fa15fac8f5cc0217fa860b60fe63f87e;
mem[899] = 144'hfdcb00ccf53df795f916f2acfb08ff38fdd3;
mem[900] = 144'h0dc4f814fc56059605cffaf707f4f4770f44;
mem[901] = 144'h08c60d7b0858faec0d85f2bdff2f0486f1bc;
mem[902] = 144'hf867044108d0fca6f49df0f404ddf8ed0f06;
mem[903] = 144'hf43008caf5080c0100ccefb0f58c0b120733;
mem[904] = 144'hfc15f90e0d9a0037eff409a60628fd8c0eea;
mem[905] = 144'hf9f8f185f85afc83f7070754f117fd620946;
mem[906] = 144'hf4a1022903fff9910775f6f80ab0ee27f42b;
mem[907] = 144'h06a8f9cb0ba6f86f051f0ef80c9bfdb2f72c;
mem[908] = 144'hf1e4f8ef0de1f969ff9bf8a3fd37faff0cae;
mem[909] = 144'hf57b0a08f1610d3d099600e303070a81f957;
mem[910] = 144'h037d0dd5024209adf5e7fa1ff78ff4a80763;
mem[911] = 144'hf376f2b305710c8af1e2ff6e030902400d99;
mem[912] = 144'h047a08aa01780819f0f305c6f11708960d63;
mem[913] = 144'hf6fafded0d1af0fd0894019301640f29fd2e;
mem[914] = 144'h0bfdfa2fffb2f621ffce04570bd8f2f70dc5;
mem[915] = 144'hf981f73f0f020fbc0656f862f097fa7cfc3d;
mem[916] = 144'hfbf4f303fe9a019e07e105fcfe660a7a0000;
mem[917] = 144'hf94ffa46fdcdff55f389f40a0d9ff765fa6b;
mem[918] = 144'h07fa01e50e6708a60c2c00fa0b6e0f4cfa16;
mem[919] = 144'hfcc8fa6004b8fdce0c5c073df67105dffd0d;
mem[920] = 144'hf71405aff5dafdd50b3deffef6cbf96f0742;
mem[921] = 144'hfcb3f5d3f1b2036af2adf6f9098e0902f353;
mem[922] = 144'hff880514f4eefab9071ef6aef916f143f77a;
mem[923] = 144'h0681fcd1021803e6f8ccf5e4f1010aeff06b;
mem[924] = 144'hfa6afe6701390d1b06e2ff730ee4f98501f1;
mem[925] = 144'h0e93fafd0ce6f550033bf442f75f09c2fece;
mem[926] = 144'hf4dc0685fc16097d09abf515f027f652fbfa;
mem[927] = 144'h06aafd9bf991011cf245f7c60214f913049e;
mem[928] = 144'hf7e3fd640f7703a403c30b7af47a083bfd32;
mem[929] = 144'hf512f9c4048d005e076cf2ea0adb0b830984;
mem[930] = 144'hf1b50bb2f9ee084e06c2fcddfacafcc00ac4;
mem[931] = 144'h081fffeaefa403f3fd42fcfc0a9e02780a31;
mem[932] = 144'h0b1bf902f823f637fb29fa5201c4f3db09b6;
mem[933] = 144'hf502fc08f191065c05dcf3c5fd5506540b5e;
mem[934] = 144'h0ec70d0003550e17f1e906be0d7a081b0271;
mem[935] = 144'hf5f2f977033cf6f906f205e2f031f6e8feee;
mem[936] = 144'hfe6807ccffcff8a6fd340b4cf5a1f2430022;
mem[937] = 144'h0168fbeaf8b102c705b80522fb18fff70926;
mem[938] = 144'hf277f7c8f1e4ffcef8e304860373fa740ee5;
mem[939] = 144'h02ea00f10d98066ffb1efc3bfbb3f9acfaa4;
mem[940] = 144'h07280bba0e62f2eff277081208ea0c5b0d3d;
mem[941] = 144'hf221fcd9f77207a7018b0a790d010f9605c1;
mem[942] = 144'h04c3fb6201240b320ed0eea2facd051ef50b;
mem[943] = 144'h0da2f754f2c0f863fda0f3d0f347fb47f58f;
mem[944] = 144'h0e170384f6a7f8c60dd5fd97fb75011106a8;
mem[945] = 144'hfcb70d3f008e04c2f6deff1a092503d3f816;
mem[946] = 144'h0b84059c058100d40741082d0e7b0bb2f0b6;
mem[947] = 144'hf9b00e83034d08160ae501ed0e41f711f686;
mem[948] = 144'h0b9af4f008b60f63f5f1f3f8fa4f05de05ec;
mem[949] = 144'h0197ff530e8d09fe09a3007907eb08460304;
mem[950] = 144'h023a0a59f7b1f3ebfa6cf00efee5f401f52b;
mem[951] = 144'h05f7f944f0e8073fff5df79e0f2402e50464;
mem[952] = 144'hfe31013ff42406280694fe05f8bef6310024;
mem[953] = 144'hf37507cd0ddbf7b804760d21f7ae0380f6e0;
mem[954] = 144'hf71cf176f8150d96f213f0b5f2abf259f21c;
mem[955] = 144'hfdf7059302cdf9f0ff940891f84f0ccdfba4;
mem[956] = 144'h06c7f77cfc60f996fdadfbc30fcc0290f0a9;
mem[957] = 144'h043cfb0eff06022c07b30a1804b90362f65c;
mem[958] = 144'hf6f80236ff9b07edfc1305b806ad0ba6fe3d;
mem[959] = 144'h03b9f38809d9009e013ff5c806d00e55fa4d;
mem[960] = 144'hffa5f8320d39fa91fa0d03c50bddf4ed0eb8;
mem[961] = 144'hf07804c8065507dcfca1f562010c0c1102cc;
mem[962] = 144'hf020f07f09d8ef8ff5d5f782f9cd0e850ed3;
mem[963] = 144'h0e5d047b093f0be0f76af2ce0c3b0baa0c57;
mem[964] = 144'hefc40716ff8cf0b1021d00e7f86b0e02f0ff;
mem[965] = 144'hf653031df46f06f2fffdffa8fcaf0082fd0d;
mem[966] = 144'hff10fb2902050503f05708c509e903ac06e0;
mem[967] = 144'hf95df75a0ec9f49701a30dcff630efaf0785;
mem[968] = 144'hfeca069ffa8101eafb0e09cc03e0f5390b27;
mem[969] = 144'hf3d9f65e0128f95400e90953014efe1bfbb8;
mem[970] = 144'hf059f8110d1af50a00fdf97cee680b180a17;
mem[971] = 144'h010af8700089f3e90350fd550853fb8e094f;
mem[972] = 144'hf6e6ffb10957fc4d06db0178f08bf48c082b;
mem[973] = 144'h027401a6fe52f9f90c77fe45f1af09990242;
mem[974] = 144'h02b3fb8afce70b9006e5fcd306830b0e03ae;
mem[975] = 144'h010807f0f1f30e95f4aff5aafe9c0126fa8e;
mem[976] = 144'hfd12ff0a050c0a7d07920263fde60da6fdb5;
mem[977] = 144'hfd5af5a0f147f877f81ffa52eff3f9ccf125;
mem[978] = 144'h067d0036059a0d9afdb3f5940d4bf058fca8;
mem[979] = 144'hfb35fbfbfc78fe7b0a00f33e07d001defe63;
mem[980] = 144'h0bd1fda603cf046af8310cb0073ffe33f36a;
mem[981] = 144'hf5baf2f6f4500d4c00c3012e085df45dffb8;
mem[982] = 144'hf35107b506a6f23af85afc93f2a9fe47f0a3;
mem[983] = 144'hfd540943f71c01210b7bf2c5fc5706240c73;
mem[984] = 144'hf537fe2e0254ff9a089b0a46037af24dfcea;
mem[985] = 144'hf1ddfd7c01020a02f807032503ce0340f361;
mem[986] = 144'hf698f9ff0a5af3caf5c90aad020b0e51fba2;
mem[987] = 144'hf61efa2af9bbf8cbfe66048a0ec4fca8005c;
mem[988] = 144'h01aa0223f1b8fe91faebf2d8f174f02e0836;
mem[989] = 144'hf011f37f0f9ff222f33e0ae70ed10757f1bf;
mem[990] = 144'hfe79fed7f674fa390b740de4f57d0ce2075e;
mem[991] = 144'hf96dff92f8e305d9f161fa69fe3ffec8096c;
mem[992] = 144'hff71f972076cfc17f6fff0b303aef64103ed;
mem[993] = 144'hef00044e0c3702fef231f2f1fb8103eb05ca;
mem[994] = 144'h05d6ff9b0d960b2fff1cf3a2f3f50d49005e;
mem[995] = 144'heeafeef60b7bf816083bece7f579092df4df;
mem[996] = 144'h09fc0547ffedf2b2fb29f7c6ef44f29b0f72;
mem[997] = 144'hf7c1f82f0659fa190bb2fc73fb3bf672fabf;
mem[998] = 144'h00ff06e7017efd9bf60cf57cf8a30499fac6;
mem[999] = 144'hf3a8f5d5f7730401efe3f302f028fe70f7d5;
mem[1000] = 144'hf942efd2f664f113019d089209cc03fd0223;
mem[1001] = 144'hf4ecf50d07770de7ef920154f8700470ef9e;
mem[1002] = 144'hff7aed2feeabfdc8edcbf5990177f1c3f761;
mem[1003] = 144'hf0f4f5f50ecbfb74ff170e140ac50388f506;
mem[1004] = 144'h0790f87ef944f353060a0ec9ff570e04f8b1;
mem[1005] = 144'hfe9b0a57f74e0c43f284f2d20e8d089b04fd;
mem[1006] = 144'hf5e2f5b6fb3afc6dedee05a9ef7b0322f5fa;
mem[1007] = 144'hfb4bf58409260d81f51bf712fc5608a60a48;
mem[1008] = 144'h014e0a3afc0ef291f3eb087efbd7f0910cca;
mem[1009] = 144'hf0f6f114056e0c6ef708fda4fdba04460a75;
mem[1010] = 144'hf504fc63046b0bd8f4810ec10d8f0d0c0757;
mem[1011] = 144'hed4afaadffacfeb4f7abfccaf94cf477f826;
mem[1012] = 144'hf2a90ef50abdfc2dfa2e00c9047af158f80d;
mem[1013] = 144'h038e088e0e2805330e3dfc80fa5bf5a3f402;
mem[1014] = 144'h062ff25afc690e2708a0054af25f0672ff73;
mem[1015] = 144'h08c0fbc70907f142f3def3effcfb064ffb62;
mem[1016] = 144'hfaccf11ffb6c0cfd0109f858f875f6ccf7e6;
mem[1017] = 144'hf5b1f8d3030ff2650287fbc1fee7f78b0d4c;
mem[1018] = 144'hff7d083cfcb40dc7ee0df5f204a9eea40805;
mem[1019] = 144'hf2b907650bde06640688f2f3f284f8550456;
mem[1020] = 144'hf363f413061f0458ff5e07fa0916003e0030;
mem[1021] = 144'h0656f565f46908c3074cfdd10aff00dbf1a7;
mem[1022] = 144'hf416f3150ae8f7d3073bf2c1f3a4f446fbb5;
mem[1023] = 144'hfda1fe05fabcf709f2290cb1f0bf09c20bc7;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule