`timescale 1ns/1ns

module wt_mem3 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h0195084a09ddf90ef089fdbf018308fcfa4d;
mem[1] = 144'h0ef50e1409220b46f45ff4d3088eeea8f760;
mem[2] = 144'h053def5e05680bf0ede2f82cfb7d0c5efbb7;
mem[3] = 144'hf8330d6c00d0090106370bcbf0ff0bdff87d;
mem[4] = 144'hf966f26bf0f2fa30030af27204bc00e1ff7e;
mem[5] = 144'hf292f6cbfc0d0df0f70beefcfbe4fb30053c;
mem[6] = 144'h0709033304fc034a040ef858f67cfa95ffea;
mem[7] = 144'hff6d02c30584ffd7f41afe39fc62f60cf991;
mem[8] = 144'h05b500cf0d1eff52000909b9fbe0f61dfc84;
mem[9] = 144'hfb82f177f0b6fbc1fa090104fa15f355fd20;
mem[10] = 144'hf066ef340448079bf09f05c9f9d3ff71f5a7;
mem[11] = 144'hfc0a0e200602f00e03e9ef350de303130b7f;
mem[12] = 144'h06ddef9e0b0d05320b8204c1f1b7ef83efb2;
mem[13] = 144'hf29a02a50ca2f111f424f301042d091bef62;
mem[14] = 144'h0e17f992005d071c09f30e040a40050f03eb;
mem[15] = 144'h074df3860666094cf93cf67af0e7f6350d13;
mem[16] = 144'hff7ff65a0e3cf04bf835f3aaf5160e7a06a7;
mem[17] = 144'h09ebfa160c9dffbff60a02dafa170d10f07f;
mem[18] = 144'hf5aefba4f430f646f2800a0cf46ef4520c9a;
mem[19] = 144'hf62cf196fa9305df0acb0ab007930bc704ac;
mem[20] = 144'h02cdf1e2f44bf5b504daf617025b02460d02;
mem[21] = 144'hfc99f43efce50f2c0f390e51fa980c20f4a7;
mem[22] = 144'hf15e0d82f5f9078301d3f994058e0ea3f301;
mem[23] = 144'hf033f5700d87fd1a0889f0b808d4f81af189;
mem[24] = 144'hfc15022f0370f0550459f616fe65ff46f3ea;
mem[25] = 144'h02020ad9fd3d09380077faabf08ef8300092;
mem[26] = 144'h01dafa5304d2f6c000b30616fb9e0398ffc2;
mem[27] = 144'hf422fddd0fbb07ca0a21f95009ef04baf450;
mem[28] = 144'hf91000a1fe07ef860424064df450fcd0043d;
mem[29] = 144'hf9de02bafd210ae2f62f0273f597ffe5fffb;
mem[30] = 144'hf5200098fd75fc2ff8c1fa48f01205130913;
mem[31] = 144'h03dbf477fe3bf3db07faf7eafd6cf617092e;
mem[32] = 144'hf49f0937ffc7fe82fd520e1ff01bf2000425;
mem[33] = 144'hf13dfaa20790f70b0595f8a5f5d1ffa8018b;
mem[34] = 144'hf3910050fa32f71df5440dfc0669ef9b0b1b;
mem[35] = 144'h0998f946f132efd804050211f8edf10206e4;
mem[36] = 144'hfa8efb3d0df304c3ff5a0af3f7b0ff2a00a3;
mem[37] = 144'h060709be09dbf19d04e1f972f78afb7afc86;
mem[38] = 144'hfe590ca4ffb9f396f065062cfda5fb8503ac;
mem[39] = 144'h0caef3650234f3d0f4a0f34cf6dbf67dfd82;
mem[40] = 144'h095c0705ff24fe79fb61ef25eefb05bff294;
mem[41] = 144'hfaf80449fcad042bf315f35bf8c7f9bb0185;
mem[42] = 144'hf3ab04d3fcfbfc80f0790bc7fcce0de6f23b;
mem[43] = 144'hfeea0368facbf950f9e8f11ffa63fe70ffd3;
mem[44] = 144'hef700618037c02a20a37091909af0782026c;
mem[45] = 144'hf3900272fbecf0eaefb901e5f806fdf604cb;
mem[46] = 144'hf60dfa50facb0ccd07cc0bddfe9bf7f9fa9c;
mem[47] = 144'h0e530dd2f34b0c5dfee3f5acfed1f4fcf78e;
mem[48] = 144'hf7a1f3e9031ff84ef1a4fe090d5009490bff;
mem[49] = 144'h0745f0eefb290b02f6c9013af45d05cbf518;
mem[50] = 144'h01ee01bd089ff38609050a8ffbbaf60efe9c;
mem[51] = 144'hfa580374fa1d0cd7f5fa058300d7ff580bc7;
mem[52] = 144'hf1450df4050e0036028101f309c5056602d8;
mem[53] = 144'h0980f561f470fe7406190a77ef8ef0ea0a5a;
mem[54] = 144'hf27ffebaf0730b57f554081900e7f6d6fce4;
mem[55] = 144'h01fbf9a205530a320891f581f6e8eff2f46d;
mem[56] = 144'h0c8b044902ff097f03faf9aaffe20c45f068;
mem[57] = 144'hfbf6056907e909f6f9fef768fb9cf7530817;
mem[58] = 144'hfeb4f6ec062f0284f692fab3fb9b09580ee1;
mem[59] = 144'hfd2301770e6f0b58f1bb052e05b90e230240;
mem[60] = 144'hf98c0358fe0dfc2efef9efa10acff901fb26;
mem[61] = 144'hf1b90a5603bb03f4fba40eb5fcf3f78cf4a1;
mem[62] = 144'hfaa2fe00fbe4069ff06e071b0154f44ff516;
mem[63] = 144'hf7e208fb0eddf68609720c5d0e35f3700993;
mem[64] = 144'h043707550aa6fbabef5af6aceef20adcffd9;
mem[65] = 144'h08d80dc40a97fcb8062504af020c075d0720;
mem[66] = 144'h0040fafa05f6f59ffa5bf14603e1f1520193;
mem[67] = 144'h0cc7f803fbe004f3fa1306de0663f20afc90;
mem[68] = 144'h0c9efe7ff1fff1550ab508170ab8f084fb99;
mem[69] = 144'h0d74f69a0c1ff4b1078ef501f43ff27c05a8;
mem[70] = 144'h05db0623f7fe0197fdfb074bf928f8d600b3;
mem[71] = 144'h0646fdb5076c0c7c0f86fed006b90790f886;
mem[72] = 144'h04dcfd95f0c30b5608d3f4e6f9380a8609e5;
mem[73] = 144'h0992f8d8028a0a96fbcbf85d0f09f0baf826;
mem[74] = 144'hfe39fc6ef66e0cea046df9fcf9d8f42b0868;
mem[75] = 144'h0e48fba1fb6af57b0e560bddf7d8f75ff520;
mem[76] = 144'h071bfa79fb2bf53406cfef260046fab2fa35;
mem[77] = 144'h003d0cbff20def1a0d63ef74f2cafa650a5e;
mem[78] = 144'h05cf0d9af56d099cfb540eb40d11fe7ff44a;
mem[79] = 144'hf61a0c3a0499f75803f10c290363f4d8f46a;
mem[80] = 144'hfff9fd9d0140efaafc6c0780f063096dfde4;
mem[81] = 144'h0215ffd1fe570803f90bfceaf463f52efb93;
mem[82] = 144'hfb660e680e10f932f78f093af9430c40047f;
mem[83] = 144'hfcaa04f609fe087df3d1f479f2ba0d49f821;
mem[84] = 144'h00ea0e98f211fb2ef7ae037d03de0429f01f;
mem[85] = 144'hefeafe1cfde2f2e50ef00ca3fda1ff500f2d;
mem[86] = 144'h0c450b7a0d90f4f3feea0dd70117f21102d7;
mem[87] = 144'hf5990cf4f84cf1d109040718fb7b0989f5d2;
mem[88] = 144'hf7ca07dc01aff1380b3f0ed50b20f24bfaa5;
mem[89] = 144'hfba4f886f06e0fe503d7ffc1fe12f3cd0235;
mem[90] = 144'h0e23fef80c8b0067006701fc089af564f8c1;
mem[91] = 144'h0ed0fb530d11004ff1cbf6abfb5df02101d0;
mem[92] = 144'hfe72fcd7f35800cff470fb3d04e607110b59;
mem[93] = 144'hf2d70d2ff8d5f4e4f90b0b08f028fbff0023;
mem[94] = 144'h0bbbfbb100260e1a02810df908d7f6240b4a;
mem[95] = 144'h04ff08d2fe6cffc0fb70f061f7ac07f70f57;
mem[96] = 144'h0ab7f8c80a0af09dfb7efe21fcdaf722f640;
mem[97] = 144'hfd07fa8ff23e0301f2bf0374f98800260433;
mem[98] = 144'hf386f2ddfa9ffc5bf0f6fc3e09f90e04f8af;
mem[99] = 144'hf2aefc37fcc8002704fe07b603200330fec3;
mem[100] = 144'hfcaefd370b3508e703dbf6bf08420c2bfccc;
mem[101] = 144'h04ed0ad50ad30181f4d3fc450862040cf33c;
mem[102] = 144'hfb140dd20da6ff390e110a710bd6fe17fcb2;
mem[103] = 144'hff9ff263f5d0074bfb5cff6f0c010da8089d;
mem[104] = 144'h0d420d170ee70febfd4d077ffcee0eec0fa3;
mem[105] = 144'hf55e0f2df614032602b402c009c807370b29;
mem[106] = 144'h0afcfa2f078df9c107b201900f0ffe0ffef1;
mem[107] = 144'h0cff0688f49e0cfe0fef011005c8002209d5;
mem[108] = 144'hf64c0dfbfdd104320e42fee3f5fe06de0902;
mem[109] = 144'hf4e7f0fcf4e60de90899f34702780e8afc4c;
mem[110] = 144'hfc3ef0f5f1970e28f87dff60f3a40733f83a;
mem[111] = 144'h0506f4b1f905fa2c01f5f741070701df03a2;
mem[112] = 144'h03610da8fd6c0e5afab90e4ffb1ff4f7ff8f;
mem[113] = 144'hf9f8f58104e8f7af09b9067100e3f6950fd2;
mem[114] = 144'hf61905ddfd1ffe15f972f084061d0fa1ff0b;
mem[115] = 144'h0a140e72046ffea90ab8f7fb03160ac2ef8b;
mem[116] = 144'hfbbcfa83f48df7660df0f80cf0f3f11a026f;
mem[117] = 144'h0ae0ff62070f055ff99e0da0fa500a70fca8;
mem[118] = 144'h082bf631075ef7da054f0e00f873fd7005c7;
mem[119] = 144'h0fa0fdaaffe8fe36f28000fff080ffe7f243;
mem[120] = 144'h0b89f29cf33afcc70423f839f733f3420f5f;
mem[121] = 144'hf1f6f2cf02e3f16ffb280e150e43ff72fe28;
mem[122] = 144'h0e5f0f38fbcc0ce6f33d0cdaf87df83a0361;
mem[123] = 144'hffd30d22f557055cf03ef4900900f99d006d;
mem[124] = 144'h093dfed8f2a00a6c0210f9bf039b0b25024c;
mem[125] = 144'h046a08adfcd5ffec023cf746f085f7d205ab;
mem[126] = 144'hfa00f51c0dcafd5a0cb7fd52f29cf1860434;
mem[127] = 144'hf0a5fee200a3f2300076ffa3f48303ddf9b8;
mem[128] = 144'hf5f8f31afccdf8040ddf0d89fc5bf7a7f229;
mem[129] = 144'h0783f239ff400a440061fa3bf03c0d9cf954;
mem[130] = 144'h018e0019fe31f047fd890e3f0144f660fb8f;
mem[131] = 144'h05a60392f9990140f3a7f9c30aff04a7fd65;
mem[132] = 144'hfc76f12df1bafef6f5c50e1908df00450863;
mem[133] = 144'h01f00c5a07eb00e4ff000bcbf132f699fe98;
mem[134] = 144'h04460f9c0131fe53fe98f9b7f1a30de1f3ac;
mem[135] = 144'hf8f0008e082cfa62fb59043d0deff9850de3;
mem[136] = 144'hfb3c0e5d05e406bc0f7503ed0fd0fc74079e;
mem[137] = 144'h07540ede0b0df4e6ffc7f8e4033d0f29015d;
mem[138] = 144'hf58d0e3e0abb09d001e4fe8afe13fc11f2b2;
mem[139] = 144'hf86a0ff5f46e0c6efb5d06500fff019b0ebd;
mem[140] = 144'hfc8c09b7f419024e06c2f015f87af72df575;
mem[141] = 144'hf9a9fe5406ba006bf285f3c8035f0db2f855;
mem[142] = 144'h04ad038e0fc8070903defd9606280ea2fff7;
mem[143] = 144'h01ea0ca301050f99f0ed0cbbff04f1eff8ac;
mem[144] = 144'h01780d5cf00f047bf78bfd440cdafb150ffa;
mem[145] = 144'hf328f1aaff510c9a0346f01709d407c3f304;
mem[146] = 144'hfdf6f0e4f9b5fa93007105ab069cf794fb1c;
mem[147] = 144'h0f760d43f43bf06807a4efc0fbbcf39f00ca;
mem[148] = 144'hf9b1066e07680d910978f1e105f4093ef724;
mem[149] = 144'hf0650398f73ff2d5f0260aea0c4f0e6809d9;
mem[150] = 144'hfc45fa70f4daf5a2fe2d077bf526f85af7b4;
mem[151] = 144'h08c50dc4fac9019f0353f11cf10401bdf20b;
mem[152] = 144'h0ae9088f0b95f90f00340c0df7bdfb2c09c1;
mem[153] = 144'hf371ff650ec103ba007708cd0c8df6790c81;
mem[154] = 144'hfcb909c1028bf884065bf2330745053309b9;
mem[155] = 144'hf491f9280990f6b6f69a0c38fb4c0361fabd;
mem[156] = 144'hf33efe4a0b2d0f11feef07370e88f402fd51;
mem[157] = 144'h07060259f6c302d7f32af5150ea80afffe7e;
mem[158] = 144'hefaa0df4f440f333eff900def14e0195f9ce;
mem[159] = 144'h057c04d00b690517fe12fa76fbba05d70fcf;
mem[160] = 144'h0bab03a4f236070a0ee7f8ccfd9f0d14f037;
mem[161] = 144'hfbf70a9f0af0fbd6f260fae6ffbdf29a0ca4;
mem[162] = 144'hf4070738ffc909cd007bf2990bfef8d4f894;
mem[163] = 144'hf8c8fac20d75f89709fcef6efd2b02c10d75;
mem[164] = 144'hf8a80ea9030d0aaff69a079804060ac0fb60;
mem[165] = 144'h06600d6df1cbfc20f1ac05e3f6330513014b;
mem[166] = 144'hfd9e009309640e9cfd54ff8a02570c35fde6;
mem[167] = 144'h084c0a84f53df6ed01780ad3fa4af2c5050b;
mem[168] = 144'h0a56058ff478f5df04ee098b0e20068f063f;
mem[169] = 144'h0ebc0c430d770d53002cfdd4f33afe96fdb4;
mem[170] = 144'h0572f1a2f968012ff0d500bc0738f927f726;
mem[171] = 144'hf0d50647f49302be0f7a04bbfa210863fca6;
mem[172] = 144'hfac10b60fc2af839f78bf9970e91faaff3f2;
mem[173] = 144'h04abfe1205160d2904f9fa940310ff6c0355;
mem[174] = 144'hf90006a4fe7cf6370776f291f4f1f6db0993;
mem[175] = 144'hf8100e79f8350e2ff26ff903f40cfc59026a;
mem[176] = 144'h09fbfbf00c65f8fb0c66f063f3bef0edfd65;
mem[177] = 144'hf28cf82ff24afb6f0761fcca01cd0a560649;
mem[178] = 144'hf49c0885ff3c086302f909e7fe54fc66075d;
mem[179] = 144'hf8470f93f341fc02f767fdc901f90acaffa1;
mem[180] = 144'hfa0ef32705810cfbfb04fc9bfb1009b908cf;
mem[181] = 144'h072bf3a90e91fa01029509c10c4603e306e1;
mem[182] = 144'h02b4ef55f1d5ef3effc0f087eff6f3f80bf1;
mem[183] = 144'hf7080a38065d0f97f158016705d6fd79f342;
mem[184] = 144'hf63eff8cf031f69403910455ff4aef190c12;
mem[185] = 144'hff430cae0ecaf64b0b49f9090806014afdd5;
mem[186] = 144'h010ff297fb66faeff101096ef82f02ee00a9;
mem[187] = 144'hf90cf3e8f43cf88f013dfb04ff7ef4e00271;
mem[188] = 144'hf73607e603f7fdd0f5ef0e3e09280b15064f;
mem[189] = 144'h000b09940eb4f768fcb5fc0df9fbf5d30d2a;
mem[190] = 144'hfc06f5d701080549ff5cf233f6faffa303c1;
mem[191] = 144'h0ee7f06900ba0c58003e04c50516f57600a3;
mem[192] = 144'hf5c3f48a0b6cf870006204eff5e908fe0885;
mem[193] = 144'hf49efe81f40c08460a8c0b40fb3207eef6ec;
mem[194] = 144'h0820f81ef9da0f09f3f0fee0f632ff87f7a6;
mem[195] = 144'hf93201d80fab0beefd1d05010c96f3d8021d;
mem[196] = 144'h0576fb83fd720c970ac6f008fd86ff2cf322;
mem[197] = 144'hfbcd09870012f34efdb4f943f64a03a4031a;
mem[198] = 144'hf8e20708f12e026df4c70ba40e97026afbe3;
mem[199] = 144'h0df1f21f0382f6b2f7a60415f226ff81fdb7;
mem[200] = 144'hfc020ce40bf0f680019c087701f8f02b0ed7;
mem[201] = 144'h0d21014c049df1a70e47f009f270f05808d5;
mem[202] = 144'h0f1ef6e60fcffe010958f2b3f0a5026b080b;
mem[203] = 144'h067bff9803d2fdb70df5f86b07effa7b042a;
mem[204] = 144'hf0c0f3830b8f02d9f3e7090d03d0fbba0da0;
mem[205] = 144'h0364fb5ef6bd093800bef2f4f55ff50af517;
mem[206] = 144'hf85cf193f876f6aa0e25f15103c5f10d0847;
mem[207] = 144'h0f0bf28b05dcf80e0d8afb43f721fd1afed2;
mem[208] = 144'h005af204f48af970082aff37f31efbf9f709;
mem[209] = 144'h0ac2f18500410f1df745fd0dfe410f6ef57a;
mem[210] = 144'hf39b0f5e074406e70dd408bef51f0c31065e;
mem[211] = 144'h045bfe620a3d0136f046f7ddfa13f666f1d6;
mem[212] = 144'hfad6f638f14df436f53b067409c2f0640510;
mem[213] = 144'h073c0c8b0e47fb42f8b7fe69f939fbcdfb05;
mem[214] = 144'hfe8af693f0e1f85401ae071c0822f7e10852;
mem[215] = 144'h0b6901d20aaef087f3c8f8e407a7fb6fffd9;
mem[216] = 144'h02f1f1ecf9ddf87f07f709fdffdbfddf0747;
mem[217] = 144'h0ed7096ffaa5f7dff750094efa0400fff972;
mem[218] = 144'h0813f2b704f0f19a04d0018105aaf91a086d;
mem[219] = 144'h07050c7605910714fa1a0138fc5204aa0ad6;
mem[220] = 144'h00c9f7cbfd09f23e0e0df1dc0be806b00e57;
mem[221] = 144'h082af2abf0cf0c42f52e0d740dba0a0cf19a;
mem[222] = 144'hf6570b8efbcb0e2f0b8702c8fb0a0c43f33f;
mem[223] = 144'hf0fc076c00a7fc41f183088bfe19017df997;
mem[224] = 144'h010f03aa0eaf0d3b053b08d20bf10794f6f0;
mem[225] = 144'hf442f81f06e4056bfe130b08f9d10b790ea6;
mem[226] = 144'hf067f2670469000cf0d4f9f605d0f3af0ddb;
mem[227] = 144'hfcd50616f0b60acb01850648f35b0c41f170;
mem[228] = 144'hf9640ba9013df843fa09f4fefbb2f3ea0ef9;
mem[229] = 144'h0ccbf6d8fae4f1d00d920c1ffa0bf8fc0106;
mem[230] = 144'h0174fb8e029905ac00670d53fb7afccb036d;
mem[231] = 144'hfa9b01e7026af111f992f7690f0509f70b98;
mem[232] = 144'hf292f6c603c80d5dfed8f7470269f1f2fbcc;
mem[233] = 144'hfcba00b706dcf8a00fbaf002f81ff3780c9f;
mem[234] = 144'hf7f1089ef846001cfbb9f45afca8f25d044d;
mem[235] = 144'hfc3ffb16fc66fc72065a038702570da00c8d;
mem[236] = 144'hfe7708ce0835f343fb64f5b9fd3f079c0236;
mem[237] = 144'h0dd30199033a09b0fd4e06a5fbd3fc970575;
mem[238] = 144'hef680de9f422f745f2a10ea7f83ffe05f9bd;
mem[239] = 144'h01e7ffedf8c10c970ded0b03041a09c6f014;
mem[240] = 144'hf6c7efd1025206de0605f168ffbbfa110342;
mem[241] = 144'hf61605dfefedf03c017cfcad0e500e260594;
mem[242] = 144'h0eb30eeef1c0fd29f37b00e2f68e0183f0c2;
mem[243] = 144'hf2c30f7bfeeaf15efc680d25fda705ab0f6b;
mem[244] = 144'hfc24fd2709e4f81c0b1ffbb2045cf1c8f57c;
mem[245] = 144'h0450fed7fb53096cf2dbfd23006e02130927;
mem[246] = 144'hf03cf3580fc4fee4fe4af26f099f05f8f4b2;
mem[247] = 144'hfa3f0d40ffa6f72b0469fcfef9e504e8fff8;
mem[248] = 144'h073bf0ce0abbf2ce040207f4fa69fb76f96d;
mem[249] = 144'hf11a0199f2f50ee40b9d0f8ef0630b65f6cf;
mem[250] = 144'h0874f3df038cf2e608b406df0d670c55f6bc;
mem[251] = 144'hfaf5099c0862f015ff970f14043cf475f26b;
mem[252] = 144'hf13ff617f1fd0888f641f7cb04cffe990074;
mem[253] = 144'hf89b07e3075ff8b6f83807b7f0710db8fe9f;
mem[254] = 144'hf461f038f9e903d008d5f6fef5510a8c0f5d;
mem[255] = 144'h0f970c97fbd6f49bf3bb0816f94cf884fead;
mem[256] = 144'hfff80a28f49efd74f9640600efff0283f238;
mem[257] = 144'h0c42f195f7c301020f140413f821fb70f181;
mem[258] = 144'hfbbc02ca0a170b91f91a08ef02da01980601;
mem[259] = 144'hf38a0f27facbf04b0a3ff7e30a52f9cef7ee;
mem[260] = 144'h0688014af99e00a5f726f258efe5f44b0e4d;
mem[261] = 144'hfdb20e560abff5c5fbeafea303df0771fb0f;
mem[262] = 144'h093df833f4f50b81f83bf539f6c60853fc0a;
mem[263] = 144'hf4dafb6b0abd0729f0acf94e0e2ff0acfeae;
mem[264] = 144'hefab05fe0f550b49098500f904d0081f05f4;
mem[265] = 144'h0ec8035b0542ff81f04f0aabfac309f70e55;
mem[266] = 144'h0006f163039c009d0b1ffcdcfb72fa420928;
mem[267] = 144'hf4d30844f722f1fc03d40cc601d8f1c1f088;
mem[268] = 144'h0b1af499ff9b0c520e050b85f05afaea0389;
mem[269] = 144'h0756fd7f04280d29fb2bfb91efe5feccf1db;
mem[270] = 144'h0b5f094cf51206740de1f4cefc96025ff89f;
mem[271] = 144'h0b18f1b00018fc73f001fb0e06b8020cfe57;
mem[272] = 144'h018406e9febd0890f7780c920091f9c9fec6;
mem[273] = 144'hfb5e08d7f008f71cf3d70a50fc820805fe0e;
mem[274] = 144'h0edc0e1409d10d5001eb0dfc04d0f5c9f884;
mem[275] = 144'h0264fa50020f065600d40439f9a3f6cafbe1;
mem[276] = 144'hf4a80005f28700f9f0a802fc0f25f08801a3;
mem[277] = 144'h01320d2af4c8f586f8c0fed2fc280cdc07ef;
mem[278] = 144'hf017f779089cf4f0fc91feb00de705d6f681;
mem[279] = 144'h09a4fd8ef6effc87f57f021e0974f537f311;
mem[280] = 144'h090ef365044cfbf8f2fa0c9900dc00480e55;
mem[281] = 144'h02d80c2a0d26f26cfbcd0f80fe2ff2b50c8a;
mem[282] = 144'hffb104ea09bcf09c0445010e0d2003030769;
mem[283] = 144'hfb99fd20f8060528078506c5010ef495f309;
mem[284] = 144'hf3390b5b0bb5f9cff2fcf6a9f3c803d50e08;
mem[285] = 144'hfd550abaf938fa2ff076f614fb2df08a0df7;
mem[286] = 144'h052505120160fc89f2cdfe020d87ef4eff7d;
mem[287] = 144'hfe3ffa1c05cefd4703c9f02c0e8709620609;
mem[288] = 144'h07e00a70fcfdf2eef0b0fdf401def043052e;
mem[289] = 144'hf5ba0b530c810b12088d045b0c56f217f462;
mem[290] = 144'hfdf9f207fa41fe3b01ecff8df4c5f6d1f8a6;
mem[291] = 144'h0d26f38cf9cefc9cf74b05eef27a00dc0dc2;
mem[292] = 144'h088c0bcff413f45b070bf17feed00b430453;
mem[293] = 144'h07f5f33ffc8c03b9f095f7c2f0f004660658;
mem[294] = 144'h0cfaf299fe4d07090154f4870dc707810b65;
mem[295] = 144'h0c6e0f3d077007020606018407b7061afa4e;
mem[296] = 144'hfd2effa8fbc403c2fb30fe3efd14f03af9d5;
mem[297] = 144'hfd20fd05fe60fd45f095f36c01a50b190a5b;
mem[298] = 144'h08c7f5510865f5110f23071309da00020b61;
mem[299] = 144'h07ccfdcbfa9af4210570f9610082089b07f3;
mem[300] = 144'h0a32f4b608bcf94af861f911f4590537fe01;
mem[301] = 144'h049706b5f395039ff375ff56f0cf07ddffb2;
mem[302] = 144'hf5d006330506f1a2f838fca1fe25fb1e0710;
mem[303] = 144'h0849025907f4fefd023d0d6404110b98f10d;
mem[304] = 144'h06dcf7b5090e04d608470eb3ef7e027e0e29;
mem[305] = 144'hfbf004c9f098f1f402ec030b0442049d0cd6;
mem[306] = 144'hf4890bd9081ef2270e220b25ff9efa1b0b01;
mem[307] = 144'h033106d900c00116fe98f2e8f83bf1490f26;
mem[308] = 144'h057ff9820b97076607e6069507b70fbe029e;
mem[309] = 144'h0017fdf9075ef401fa5d07b1f67809ac0e34;
mem[310] = 144'hf7bdfe12065bf010012803f1f4cbf0fbf582;
mem[311] = 144'hf3fdefac0764f104f784036a00acf0d703d1;
mem[312] = 144'h0cc1fc7206dbf9d8fbda042ff0bb04230f77;
mem[313] = 144'hf1a5014a063ef9b00b6ff279f66df881fb3c;
mem[314] = 144'hf1ff0e7a02820d0c0bba0b92fa450a9603cb;
mem[315] = 144'h02180bb207f0f5f5f6b6fcaf0de1012df3d9;
mem[316] = 144'h0a89f7baf7adfcf1ffedf779075403d9fc9e;
mem[317] = 144'hfae6fe90f27ffef5fb4b0430f997f2ae0964;
mem[318] = 144'h0083f55ef854000e0468f955f8b405cdfdab;
mem[319] = 144'h0ee5fd15f7a80fc7f552f157f35b01f50729;
mem[320] = 144'h0a4b0b2e0a9cf9b907320fa8f9b2feaefb53;
mem[321] = 144'hf8230a390144fe94fe480b070bd0f02701ad;
mem[322] = 144'h0cf80be8f780f0fcfd67f6ddf4c507dff629;
mem[323] = 144'h04bf0b4bf713fa7eee9e08600cc4f2ca0482;
mem[324] = 144'hff6ef072f3bbf30df07afeb50361f538f98b;
mem[325] = 144'h01360c1a03edf5fe0cd9fe9309e3ef0a0c32;
mem[326] = 144'h042404700899f249f0c1f99af0d604a608e0;
mem[327] = 144'h0a7cfe2d007e048604ef0d6703cbf121f510;
mem[328] = 144'h02100e3b0475eef6f51df52502d607660247;
mem[329] = 144'hf87df92c0f6507650334fcd9f85cf169f946;
mem[330] = 144'h06d30d50f0e60ec708e406b50ac2f3e9fd90;
mem[331] = 144'h01fb03cf00e5f3390ae6f5fc0bae0570085f;
mem[332] = 144'h0cf305a00f1e010601e6ff86089e0949ff1a;
mem[333] = 144'hfb07012a099404d2f61afd69f4a70750fb16;
mem[334] = 144'h01460d8ffac10978feb1fb4508ce08770ad5;
mem[335] = 144'h069f07c9007002a90e9ff873fd2109c40ca6;
mem[336] = 144'hf8bf0f17022cfe3a0b32013a04fef185fd64;
mem[337] = 144'h05fcf1310ba605a8085ffa04014bf41900eb;
mem[338] = 144'h03cf019cfec0f1f4f503f54309fafc000e16;
mem[339] = 144'h0dfbfa6505360d62088df9fe0de0f7d40855;
mem[340] = 144'h08a70a0b04740d760f1df77bf0e5fb6c0b7b;
mem[341] = 144'h02530e0909f50e68f14c0400f614081bfa6e;
mem[342] = 144'hf06d0fb8f052f0c2084e0a9d0e07f5edfb37;
mem[343] = 144'hf8c6fc77f5b60389fcf9fb0aff3a0ad60c8b;
mem[344] = 144'hf640fa2cf6090771f26af20df3cffdbe0921;
mem[345] = 144'h0b61ff3af8c401c2ff4103b1f1f20f87f44b;
mem[346] = 144'h08d40eecf1cff96ff7be0c2ffff40e3f0b8d;
mem[347] = 144'h069ef1090719f46ef938f9e1077801e2f2a1;
mem[348] = 144'h08d1039c08dff4030a7e0cc7096ef4490e6e;
mem[349] = 144'h0e17feb007a508f6fdcf0d3607580938febd;
mem[350] = 144'h0779f3daf8230be00cdff7bff059f7b10a61;
mem[351] = 144'h06e2f3950a450cc2fb6f0e2e0c61f6c7fe5a;
mem[352] = 144'h0197f138f7dbfc120e1d035b07450cf6f31e;
mem[353] = 144'hfab2fe89f872fd2d0c18fc61f4770c130197;
mem[354] = 144'h01eefab8fe030b23f334018afd36f47e0965;
mem[355] = 144'h00c00d35faf5f779f52500ba0393026cf3b2;
mem[356] = 144'h0260f174fd8008cd0dca0644f2d9f861ff5f;
mem[357] = 144'h00f00d8bff7ffc32f4a7fccbf84ef35af7b3;
mem[358] = 144'hfcbb04e90e580a82f2480aad04f4f8c7fc7d;
mem[359] = 144'h0e1ffdabfc3a0f7803c20425ff0afc4ff087;
mem[360] = 144'h050afcfcfbd0f0800153f5aaf050090f010c;
mem[361] = 144'h04d7048bff4afff2fb2ef4da0487fa3bf221;
mem[362] = 144'h0ca501f102c2f52cfa6606d1f08303520bd0;
mem[363] = 144'h006af6daf30b0b17f1d70d2f0f77f8860416;
mem[364] = 144'hfc43f00806b70ec90b010141facbf2880cc1;
mem[365] = 144'h0014fc98f04208ee0c040e7cfec60d46f5a1;
mem[366] = 144'h061f0ebdfac80aedf71ff3d40936025dfe49;
mem[367] = 144'hf03a0a25f7a7060af8f3fca700f7f517f53f;
mem[368] = 144'hf722084b0c7c0b17064a05850be60739f728;
mem[369] = 144'h068ff2dd097af619f9f403020615f865047b;
mem[370] = 144'hf44408f2092109e5f6a3fbad05d209f50be8;
mem[371] = 144'hfa8900e0033d090e0aa10d3ef211f209f84d;
mem[372] = 144'hfdbf070af654042a021c0c7f03c70c860e54;
mem[373] = 144'hfc910f8bf14b06c101240b37f2fd01df0e0c;
mem[374] = 144'hf9e5037b0060f26ef0cc034efe990627f411;
mem[375] = 144'h0772094d001b0a78081cff24f9ff0a43f380;
mem[376] = 144'h019c0d21f2fb0b61f68beff7f87aff99f485;
mem[377] = 144'hf7b6f8fb02220100fdc4f03bfc29fc050731;
mem[378] = 144'hf25ef7d10258033ff563f6b5086ff66ffe1b;
mem[379] = 144'hf8750b03010106b7049e0b2dfd570b0df36c;
mem[380] = 144'h0f05099509bbf0230a9bf080f56af57c033f;
mem[381] = 144'hf86ff7ce0beff7880754f74006eb01a0f628;
mem[382] = 144'hfc9bf9a2f5d5fe02f0c305a9f3ccf584fd6f;
mem[383] = 144'hf218060df30e0ef50b8f0aebfcb0fc8a0b42;
mem[384] = 144'h0628f98805f50bfcf4c007f40f0a075e0756;
mem[385] = 144'hf2610201f771f143f31bfc58f89df6e6fcb5;
mem[386] = 144'h0adefb8af8f906caf48b091004fe01050a98;
mem[387] = 144'h0e270113f129fcc0fe55f43cfd7d0e55f108;
mem[388] = 144'h007d0d500184fc2dffcbf0a60b970669fe60;
mem[389] = 144'hfd670f250ec80dbb0421f6bc07b607d00237;
mem[390] = 144'hf4eefe8c0b54092809aaf110f5cff1f6fac0;
mem[391] = 144'h0d5f0e920494ff4bf77d07c2f58bf614f5b7;
mem[392] = 144'hfde5008d08b0f676f06cfa4a0d0b099bf3b9;
mem[393] = 144'h06500e98fb81fc4501ad056af7a1052a0489;
mem[394] = 144'h0663fc1a0988f135015e03c607b60730feeb;
mem[395] = 144'h054b0ae9f682fc13089c057f003cf7d9fa52;
mem[396] = 144'hf0b80eedf3700e8efe16f841ff740eeaf810;
mem[397] = 144'hf845f40e0cfffab4efdcfad00560f6ab033f;
mem[398] = 144'h07c4f029fdb8f35f0934ff17036606a7f4a1;
mem[399] = 144'hf71b0838f03cfaa5f8d1044a07ebf616f184;
mem[400] = 144'hf4b2ff1ef2b0fbb40b39fdf6f3b2072ffcb9;
mem[401] = 144'h0b5e0132fd28f255fb59011bf2c0ffcaf703;
mem[402] = 144'h004600710eb20191fc17003bf1cf0a66022c;
mem[403] = 144'hf7d5fd29fd2cf859079e0b06ff88fce8f49e;
mem[404] = 144'h0366fc4c0b25f89ffdde039904aafc5507df;
mem[405] = 144'hf127ff23f95e0c6d0a340d88f145f212048f;
mem[406] = 144'hf71cf9560eee0902f4d20d410685f912031b;
mem[407] = 144'h099a07730645ffa4f29efe1300630066f96b;
mem[408] = 144'hf32d0064eff80671038e0dc8f2bf0b67ff5f;
mem[409] = 144'h0ca005e0f6820b2b071e092cf32a082df270;
mem[410] = 144'h0075f817050afe5ff816ff44079f0d96f9c2;
mem[411] = 144'hf606f472f122f1c405160a480a59f6800463;
mem[412] = 144'hf020f9180892f21ffaa50d6ff3550a380834;
mem[413] = 144'h0870f86cf78201a7f3c8060ff4150ae8f946;
mem[414] = 144'h0cc1fca6052bf179fc9ff3c9f593fe96058a;
mem[415] = 144'hfefb07be00e60361fc45ff2efb4101ad0304;
mem[416] = 144'h0ec6f5dbf498f0500ac2f4bdfd0bffcdfca2;
mem[417] = 144'hf351fc98014f0c150586fde30522fe730af2;
mem[418] = 144'hf164f280f2a9fff20ad70aa0078bf4d4f797;
mem[419] = 144'hfe28ff13f17402ecf168088bfc6b092a0311;
mem[420] = 144'hf3b708f6034b02f9ff1d0f020559f672fa79;
mem[421] = 144'h0448f3a6f9deff6bfeeeff62f11bf8a70843;
mem[422] = 144'hf9340287f30b029bf31fefbe044ff498ff26;
mem[423] = 144'hfe67f087f9770f40f1ccf971f279ff17febb;
mem[424] = 144'h067c023f01480390f30e0836020b03cb0859;
mem[425] = 144'h0e2af4c4f251f66f08c7fcf80d6709a80aa6;
mem[426] = 144'hf3dd0e280c13f16803c102a9081d0e53f04a;
mem[427] = 144'hf88c064df155f2c4fd2b077d0056f2a5f87d;
mem[428] = 144'hf25f000609940347fa5f0ef6f26ff59bf532;
mem[429] = 144'hf683f138f0d902cdf7e00c38084e0690ff78;
mem[430] = 144'hf7dbf3870e00f8760427f27705680a8ef283;
mem[431] = 144'hfc9c030f0b5d053ff6340b940419099ef749;
mem[432] = 144'hff9fffacfa96ffd8072cfcd2feae0be40a61;
mem[433] = 144'hf7aff413fb0c0394f5d80b16f3760a360f40;
mem[434] = 144'hfe2afef80087f5f5f44c032df8dcfd5703f2;
mem[435] = 144'h0285022d0242027a07eff015f7e70ca7f5c7;
mem[436] = 144'h01bff4290de20c84fc06fd67fb14f894fa8a;
mem[437] = 144'hfb55f96b0dba0c5df2dd090e016af3d1f56b;
mem[438] = 144'heefe04fb026bf70af436feeefe91efb700ee;
mem[439] = 144'hf166ef35ff4202230a3cfc00f934f8e0fb7b;
mem[440] = 144'h011efe3003eef596faed0cd1f7180f1b0625;
mem[441] = 144'hf343fbdb0475fd10f865f4640989f7f2f477;
mem[442] = 144'hf14cf6720d2cfe6e0cc40a3dfb9af6b9ff1f;
mem[443] = 144'hfacff8380d7afbcff9dbf2bd06e0f738095d;
mem[444] = 144'h007607d4068af939f5c2050cf4ca0560f183;
mem[445] = 144'h0e070480079ffe4702960ec0f0eaf91a0c7f;
mem[446] = 144'h0478047d05a7f748f144f490f224f125fd58;
mem[447] = 144'hf287f5adfd9ef8660fb9f045f3bb0a81f87e;
mem[448] = 144'h013c05dc0773f379ff01f2c5f42ffa54029d;
mem[449] = 144'hf36c09def21d0b17feecfb3df427f5d5f0a2;
mem[450] = 144'hf9d20462049308f7f9c30e2efb06f35efd26;
mem[451] = 144'hfebfeffa021ff379fe07058cf984037b0725;
mem[452] = 144'h034e0101079e04abf9bb0fb6efe6043b0407;
mem[453] = 144'h02c3f10a0cfdf2e6fe22004af00e0e09fa5b;
mem[454] = 144'h089005c4f2d0f14df9fe03e5f653f09c0c89;
mem[455] = 144'h02c8f0e50c8d016efe74f832ffb3fa1df486;
mem[456] = 144'h0d8508bafef2f3da02b306ef02d9f736f170;
mem[457] = 144'hfcb6f9c3f365f81e036afc970001fc05f736;
mem[458] = 144'h0c4f0c26024bf00a080c0cbeffd408b6ff72;
mem[459] = 144'h0752f77d0343fa1006eaf2850e6b0f410330;
mem[460] = 144'hf066f5da01c7f655f596fe0f0062f33c0170;
mem[461] = 144'h00d6fe7d0a2f0ab5f31ff126f2e1f9fefcf4;
mem[462] = 144'hf853f20803a904eb0c4af6c20398fbf4fafe;
mem[463] = 144'h0bdff9bf0c670c16f5f802f1fea80e130d13;
mem[464] = 144'hf705fbb9fb670225f3ef0b3df822f2ea0e1d;
mem[465] = 144'hffd6048708890f420258fd9300ceefc0fe72;
mem[466] = 144'hf337f833f3e1f4c0ff120695fdcbf4ae033c;
mem[467] = 144'h0d99072c05850e8708e2ff1f02b6f322f83b;
mem[468] = 144'h02bff6aefeae01500c1fffb50a4904690747;
mem[469] = 144'hf4cd0f650c000556f31109460903f0ebfbeb;
mem[470] = 144'h0a3cf9c4fea401340a3701480a0608a2ff5e;
mem[471] = 144'hfc93f83afb4a04a5fe13fe860c2c08aff3e5;
mem[472] = 144'hf6dbf7cdf25d0492f5d40640f70def97fad3;
mem[473] = 144'hf977f1ad0d4e0149f3250016f394f55d05dc;
mem[474] = 144'h0065fc390b05f1790d6ff5240910f96802c5;
mem[475] = 144'hf99a02e50395f7cdfd7cf425f1cff569f5c9;
mem[476] = 144'hf9f5030507cd09fcf9e2f0710a6af04d0ed5;
mem[477] = 144'h048bfe47fe2ff3a9fa98fdeffc1bf8f4f8ca;
mem[478] = 144'hfbda05fb020bf6340ee5f650027901e8f71a;
mem[479] = 144'hfdea0d6c0f1201e004190a5e0342fae1f563;
mem[480] = 144'h05a10071effdfb6002ed053702a9fa930666;
mem[481] = 144'hf871ff86078ef4830b20fa34f9060c07fa96;
mem[482] = 144'h009dff5df667f903f48f0f360942f61c03d7;
mem[483] = 144'h0716fcebf505fd01fe62f783f986f4080403;
mem[484] = 144'h06b20db40557060a0b9ef1580cea0720019b;
mem[485] = 144'hf819ff44fa38f7a70c2bf65c00480c15fc6e;
mem[486] = 144'hf7300a8c0cbef175076f090afc450b81f43c;
mem[487] = 144'hf59a0f6d004d0536f6e5f02307acfd43fef6;
mem[488] = 144'hf6b407db027e070302aaff5cf7ae0641f771;
mem[489] = 144'hfe7c066ffa5d08aef2e702ddf7e00c39f770;
mem[490] = 144'hf990f6c1fac90e4d0fdff70bf21c09c8f6da;
mem[491] = 144'h0c6d0dd00ad3f8b60819fdc0098cf658f711;
mem[492] = 144'h05b3f807038c09acf3960f350c4eff67fc30;
mem[493] = 144'hfe2b02edf32df2f6034eef85f20608a5f1ed;
mem[494] = 144'h0e5f0e75fb15f8e104e3f5bafed807a7f44b;
mem[495] = 144'hfed2ff82f2bb0ac106a5038107220751f9de;
mem[496] = 144'h0e97f0b3fe35fd06f3cc0f7a0c7902e0f592;
mem[497] = 144'h01e2079d074cf0970baf0dc4f4b1f937fda8;
mem[498] = 144'hff3c0b69fcb3f5f70937f9f30b3cf266025c;
mem[499] = 144'h0b65087d085d052702ce0ccdfb0af272f63f;
mem[500] = 144'hf1b8f366f2c7f0cbf8b2045ff1250dc0f099;
mem[501] = 144'h050f0298fbcf0933f045feed0b2609bb0250;
mem[502] = 144'h0332067df4500092fb55f6aa05acfe47fc29;
mem[503] = 144'hf96df002f78302f10190085cfbd0efb902b5;
mem[504] = 144'hf3c4fc010bae0ddd09220cd2065f0470fc52;
mem[505] = 144'hf674f6c20b39f805f3510170f248f93a0301;
mem[506] = 144'hf8ff0ba7037dfa8ef161f72d056d0d30f122;
mem[507] = 144'h071806fdf381f69e0d73f3c5f7a1f132f7bb;
mem[508] = 144'hf59b096cfae003ae0d13f7fe0d78fb87fc98;
mem[509] = 144'h0c5b0c00f0a403d8fa2b0619fa2407240671;
mem[510] = 144'heee10792f4e40511f0d6fee0f8db07290bdb;
mem[511] = 144'hf82afef10f96f7f4f8a4f9d5f2ad09490a29;
mem[512] = 144'h0da3ff11f22301010667fd0f0f2000ca09fc;
mem[513] = 144'hf644f6af0a85fd23fbe50100ef5ff3fef61f;
mem[514] = 144'h06750ba5fcec036df267f8f80b0a0b80053c;
mem[515] = 144'h0a31fe51ffc400ddf725fbfafc8b0abef468;
mem[516] = 144'hf2b30ab5f420f3fb06b3f8cd0965fb89f809;
mem[517] = 144'h0892f4f2fe27fe8af15afcbef3310041013a;
mem[518] = 144'hf9f704650a0702c1fcb60854f35207ca0aab;
mem[519] = 144'h0d6e01e4ffc3070f041806a5f6abf7210aaf;
mem[520] = 144'h08dbf813f4f70ca50d4a0d9a0345016cfdee;
mem[521] = 144'h04dcf9790265f9b4fae70ea9082cfccffec5;
mem[522] = 144'h0aabf08e05dcf904f55f0f9df0d3f7b30a0c;
mem[523] = 144'hf183fa62f2040df7f628018cf9a6002cf079;
mem[524] = 144'h0208093ff5af0389f71b0e8df552f9c8f6c0;
mem[525] = 144'h0ad9f9110a03f3950895f052f4e2081502c3;
mem[526] = 144'h07470d950a260a8af239f98cf4bc05480038;
mem[527] = 144'h0e9605380965f20bfc6dfd85f1d8fa3f0720;
mem[528] = 144'h095b093b07b5f527f7ae0c1efbdefbbe076f;
mem[529] = 144'h0bf60b8cf1f80f94fde1ff5006e9f53109df;
mem[530] = 144'hf4bc0e86f57a0238fe84f81e0c90ff6400a8;
mem[531] = 144'h0cdc0d360ab7074401a60ad5f7c80c2a06f4;
mem[532] = 144'hfdcc0af4f95706f9f88a00b3ffb40a00f58a;
mem[533] = 144'h0b430163f79b03c0efde037c0a6a0c1d065b;
mem[534] = 144'hf3bb031d0739f97dfd4bfd530d3507010d6a;
mem[535] = 144'hfd8ef112f5eaf2b5065b0e1607250c43fcb5;
mem[536] = 144'hf997fee80391fc05f501f20308290ea5f43b;
mem[537] = 144'hf17e039ef96a0d55fdd8f92003b7fb03f39d;
mem[538] = 144'h04cef7940bd0f60c0bfc0010f48b0dfdfaaa;
mem[539] = 144'h0bd8ffd7f39d0e0c09e50ea40c5c0906071f;
mem[540] = 144'hffbc0b9ff39e014d0110fdf70902fc20f886;
mem[541] = 144'h0bb8f826f2680bdd0e10027f043d05e00ec0;
mem[542] = 144'h0a59f77cf094ffaffef40b53f1860e0505c6;
mem[543] = 144'h0bc90a6608ef08a102b3f61d0a57f8b3f24b;
mem[544] = 144'h0e690f5af53bf7e50eaa061b0d9008290085;
mem[545] = 144'hf7c4f6480f3df1960a49fed8f03def2afeb8;
mem[546] = 144'h08ea027af7a1099a0d1e0504f8190bc2fb30;
mem[547] = 144'h0661003ff932050df94a0a550b90fa01f905;
mem[548] = 144'h068b0bbe0dd8fcd40f55f83bf8dffd7ff746;
mem[549] = 144'h0a47fc0cfb820b40f9fb078e0850f7eff8c7;
mem[550] = 144'hfb0706d4fd2cfba4f7fd08fd012bffd60820;
mem[551] = 144'hf7e20051f92702f0f770f389f77602c70165;
mem[552] = 144'h04e30230079bfd89f5d0012d035bff79030b;
mem[553] = 144'hfdbff24dfa87fa8f0df1fb5afde303bef9d3;
mem[554] = 144'h03da05ae0e5707b9fc44f0bf07d90dcc01ca;
mem[555] = 144'h036ef9a50d6d011df5bbf500f2aa00390002;
mem[556] = 144'hff0c0757f29a06ac09d7f5f203420ad90dce;
mem[557] = 144'h0b2ff4a601fbf52a0155fde9f74b0003ffdd;
mem[558] = 144'hf752f4f200a60ac1f9d30a35f143f3c4070f;
mem[559] = 144'hf365fa0c0c9ff9e30be0f292097f0f9afc7b;
mem[560] = 144'hf8b506d70b520eacf54dfca9fb2a0322f49f;
mem[561] = 144'h08360b67f4d90ed608070d62fa26033f003f;
mem[562] = 144'hf2e90754fc7400160f2af8870a74fe100cdf;
mem[563] = 144'h0d8a00b0049a022408b9064bfcfff51cff31;
mem[564] = 144'hf2a102600fb0f21a0d9d05d30e890118f634;
mem[565] = 144'hf6e3f21efe3dfc69f7e4f7a7f110f8640da8;
mem[566] = 144'hf668f625f447ffd3f165f1d3f8ae09eefdd1;
mem[567] = 144'h09f900e5fca4009bf75b0e540850fe1cf68a;
mem[568] = 144'hf8e50f36f78cf7eef424089af1dc0b44fbdb;
mem[569] = 144'hf55cfbccfefc012c0c8f06a0fc09f6ae030e;
mem[570] = 144'h09f705a9f2ecf69cfb8502b3008801c00a6d;
mem[571] = 144'h07210769fb5ef69905e2fe2bf84afe040aca;
mem[572] = 144'hf02cf15bf3780564f596f99e0806f21a04eb;
mem[573] = 144'hf7d5feaf0da104eb0831f2930c420099f938;
mem[574] = 144'hfd6d07730b35038706010470f63dfb60ffd3;
mem[575] = 144'h06520e2ef7d6092dfe97f744f8def2c2f2f2;
mem[576] = 144'hf25304f6f2aff27d06ae0adc0af8fcb0f0bf;
mem[577] = 144'h06c1f51bf441f41706abff49f8db0996f53d;
mem[578] = 144'h02430ea509c6f88507acfb32f4ab02fe0871;
mem[579] = 144'h07be0ca0012b019407fe0a29029dfb2ffe94;
mem[580] = 144'h01e0ff680e08f21802e3f1f80a59f7dffa45;
mem[581] = 144'h057a08200387f132f338f4b1f059013d0a5e;
mem[582] = 144'hfedc0f410badfdcb0ea00641fd7709e7f160;
mem[583] = 144'h022bfe5b0f91f3e9f9edf6c20e930e22f67a;
mem[584] = 144'h0d1afe63f312f126002c076d0ee1f9db079b;
mem[585] = 144'h054d041ef8260c37f6fb04830a43fabcf595;
mem[586] = 144'h08c2fdccefe3018dfbb2fe80f728fb7e0854;
mem[587] = 144'hf973f55b0e73012f0bd2fd9a075b0a710bda;
mem[588] = 144'hf1e3034aefaf0ea006b2fe9ef26b091dfe35;
mem[589] = 144'hef030ba108c8fde0f68ff137083af297fd4e;
mem[590] = 144'hf4fffb0afa660d89f9760c95fd6c0ed40c42;
mem[591] = 144'hfa4c07c3f373073007eaf08c00390c90f974;
mem[592] = 144'hf5330ac7f00c004506af0613f04ef486fdcf;
mem[593] = 144'h0b75f4bf0e5bf8cafac0fbe9f6cf0e3a0442;
mem[594] = 144'h034afa75f98df393f362f23ff0680aef08aa;
mem[595] = 144'hf5c808e408300d790f94061efa45fdf0f913;
mem[596] = 144'hfff6078b07e9f5000cd1fe4ef8b0015afe87;
mem[597] = 144'h0da90c1c0236fd030b97f49306d7f2650292;
mem[598] = 144'h063608d50ba705fff1400c4af5e607a70ac2;
mem[599] = 144'h04a40540f0ce0254017106a0fa250441061d;
mem[600] = 144'hfb7d07250eee007df6aff84cf5680c51f53f;
mem[601] = 144'hf8210a2af485fe4402bcf7920803070d0bcd;
mem[602] = 144'h0d1df7d2ff39f70307ed0684f95ceff6f2ce;
mem[603] = 144'h0e8f0359fd410dfa0ab800800671f12e03d7;
mem[604] = 144'h02dbf2de0c8f0be5ef6a05830aa402d1f5a8;
mem[605] = 144'h0926fe93fa640054fcac0303f2170cadf94c;
mem[606] = 144'h01ad0288f5a40d6e097eff870e3a05880afe;
mem[607] = 144'h0ff409750f77f2a30ddb06bd0070f328f6e8;
mem[608] = 144'h02a3034bf9e5090df3dc044a009403ca058d;
mem[609] = 144'h05e2018a0b7305560aaef63b0ae0048a0228;
mem[610] = 144'hfc24f63a0bb1f241f2930efff4b70bc2fe4c;
mem[611] = 144'hff7afc41f3dafcee09a8fd7b0dde0985f142;
mem[612] = 144'h0bb3f8bff7330675faa9018ff145f99bfab0;
mem[613] = 144'hf007fefdfb52f5700a4f048ffe800661f10d;
mem[614] = 144'h023004d2013ff94dfd570c130be30709f442;
mem[615] = 144'hffbef02af8d2f2850518f6420414050bf39a;
mem[616] = 144'hf54ffbce05b70bbc0c3afa04028400e00515;
mem[617] = 144'hf0680ee2fc37f6dc0ebb07f907e7f062f396;
mem[618] = 144'hf5d50a07f5dd08cbf27bf5d4fc03f9bdfa6b;
mem[619] = 144'h0d0600d0f68bfce2f5fafd34f1f80db1f2fc;
mem[620] = 144'h0479f81a06cffd2ef89c0ec2f396f1f10805;
mem[621] = 144'hf053f8d10c78fb940307fed9fca7fab9ef74;
mem[622] = 144'h0adb0dc10ae0f3fc03ecf4fb0cad061603ad;
mem[623] = 144'h0d1cfa33f61cf2dc0bd2fa45f378042cfba5;
mem[624] = 144'hfd7cfec5040a0c9b083c0c360ca7f952f6f4;
mem[625] = 144'h0937f667ff90f002ff110a610d76f687056c;
mem[626] = 144'h05a5f9450a2308620cd4086e08f50b8affec;
mem[627] = 144'hf1a2fbe4f0b6f82e04050d06fa830dc9f85b;
mem[628] = 144'hfcb2fa5cffcaf6d908a7f41bf41c059efa66;
mem[629] = 144'hef21f988f377fe38f3a207b4f988fc25f68a;
mem[630] = 144'h00fbef480d65fb8302350cdf00f6054bfe22;
mem[631] = 144'h04f6fe94fb56f841f789fcf9f544f13df2b5;
mem[632] = 144'hf9c4fdc9fa92f104efe8f7db027afddff02a;
mem[633] = 144'h0b9b0a55f18dfbccf074f9e30c52f663ff1f;
mem[634] = 144'h02dcf8a7f098fa3ff44b0bc1f4c0f70704ff;
mem[635] = 144'hf9040c8a05f00e2f0a6009a80213046fffb7;
mem[636] = 144'h0840f953f0ca03410739fa5eff3bf2b9f76f;
mem[637] = 144'h0097006ff26b08d8f9d5ff2f05c2044b0339;
mem[638] = 144'hf3d5f1bd0d1e05fef602fe890966f3c70da2;
mem[639] = 144'hf33f09e005250e910908ff11f9f8fe77f41f;
mem[640] = 144'hf9cef2eaf12507defeacf9ccf4c9f6230061;
mem[641] = 144'h0d83f0cc0743fde704da05b408f504a9f552;
mem[642] = 144'h0d100c7c07950e15fb92fcac0d9000b1fa2a;
mem[643] = 144'h04d204d808320181f0fff681fa84f7ca0c67;
mem[644] = 144'h0d95f2070e280335f8a90735f7820051fe5f;
mem[645] = 144'hf4ccf4d0f4e6f89ffa03f9aefa6efc210798;
mem[646] = 144'hf9f5fa66f5d108fcf1eefe36fca0023b0833;
mem[647] = 144'hf1cef143f35e0c1e0f500e63085200600d3e;
mem[648] = 144'h0bb40acb0452f69df23aff46f984f8940503;
mem[649] = 144'h0fc7047e0f1f00bd08de03e2f125ff70f11e;
mem[650] = 144'hf32bf6ea0d21f420f27b003dfc61f2250a19;
mem[651] = 144'h09dbf0770003f7010972f9fbf21af1cd0c60;
mem[652] = 144'hf1530d1d0f180a0c068cfd41023601aff352;
mem[653] = 144'hf46e0bb30ad1f006fddbf6600de3f7a7082e;
mem[654] = 144'hf07e0329077bffdb01d5fc880c23f23cface;
mem[655] = 144'h08910e8e022af0ecf526f7ccf9090dd404fd;
mem[656] = 144'h002e07f50d420a860c30fea2f7e40ba4fd08;
mem[657] = 144'h0896f7e00b1df79b02e4f2df0aa60b5a0d91;
mem[658] = 144'hf1ebf616f301f2a705480e9e0bc4f79bf8f1;
mem[659] = 144'h03b30cd404a3f7c0faf802d7f580f779f88d;
mem[660] = 144'hffcb02e000650ebdef7fff51f5ee0c31fe9a;
mem[661] = 144'h0c7deff309c1fc36f7bf01670ee10ee6036c;
mem[662] = 144'h0c6f0b5a039df434fd8608d0fd2b0d7f07ef;
mem[663] = 144'hfe97f558f6aff470f50d0760ffe6091c06fe;
mem[664] = 144'hf24805cc03a7ffbffbc9fb7cf9ccfcf5fd39;
mem[665] = 144'h0d8707780efc0846f2f0f930014e01000d6a;
mem[666] = 144'h0ca400f10e87054503950daaf35f00a201bb;
mem[667] = 144'hf3ca0176f907f539f2fff111f753f3340023;
mem[668] = 144'hfb06ffe4fd040665f18f0a960dd7f9ed0226;
mem[669] = 144'hfee8fff4f59d0c55f360f20c09390e700d24;
mem[670] = 144'hf4acf3e4f2000420f20cefe60d280dc30e3e;
mem[671] = 144'hf03203ca0f13f1a20ef5035a034ef2fcf991;
mem[672] = 144'h0833ff66fa9d01abf7ecfcf8fc630c24f12b;
mem[673] = 144'h0cfafb150891087df0dc009d03ecf0d3f729;
mem[674] = 144'hf7d006100bd8098708260a09fc38f8070c24;
mem[675] = 144'h0933f928068803f005fbefe5090cfef40944;
mem[676] = 144'hf59af4e70da1f1630503f64efc20fb4e0cf7;
mem[677] = 144'h051bf2cb05bbf8160bfb0eb00b81f0fd00fb;
mem[678] = 144'hf224f2690074f525fbef04330e86ffe9fbf9;
mem[679] = 144'hf76f093805b7fce6067ef5ec02b900bf08f8;
mem[680] = 144'hff9d04dbf262f1a3f7d808480aa9fbd9efca;
mem[681] = 144'hf04b0aae03b6f5b1fb5cf980f4a70d810bb0;
mem[682] = 144'hfed703a3f60f0ec301dafae80d18f491f179;
mem[683] = 144'hf729044efab7f4c9060dfc04f23e096b0b8f;
mem[684] = 144'hf7daf757f806f595fc7ffc8704d3fcd0fb3d;
mem[685] = 144'h0052f5cb0702f0070bfdf7bc0da0ff940746;
mem[686] = 144'h07eb01600855f2c50cf90d850833fbaf0552;
mem[687] = 144'hf73e0944f8f6073ef243f1960d77f990f14c;
mem[688] = 144'h0086fc010ba60c8cf0970a980d96fcfbf4ea;
mem[689] = 144'h0053f0b5fcdd030d00a7f3cd0d5cfe570922;
mem[690] = 144'h0a820e40f4cc0fdcfa8b09e9066af1c2f617;
mem[691] = 144'hf69efb76f6e806d207cd03a7f941f74e08a8;
mem[692] = 144'hf7c4091e01350cfd00910b610e08f1d50f02;
mem[693] = 144'hf6b1093df7e70ed3f4c4fba10f61f41ef3a2;
mem[694] = 144'hfbd404640dbcffab05de0a54f3a0f3360ff4;
mem[695] = 144'hfcfb0f67f4470f62f46df5ca0ec201b60b20;
mem[696] = 144'h06ac08030f52f537f62afc7807e3fe3a0167;
mem[697] = 144'hf1aa0b03f79009cafc48fdf8f5fb08be0b57;
mem[698] = 144'h080a07b001d00dc60a2006bdfc01fc1f06a5;
mem[699] = 144'h06ecf5510e66f463f23608840c7afb07f63e;
mem[700] = 144'hfe14f434fd1300d10fdd0a5cf163fb5ff1e6;
mem[701] = 144'h03330b1104a7f11cfdef03540fde0b570704;
mem[702] = 144'h0c43027e005bfc48f094041af892022a02d9;
mem[703] = 144'h049cf9d0f43cf72e027904e90e4c0cf0fed9;
mem[704] = 144'h08a0f00cf8560821ffc101a8f695f473fe83;
mem[705] = 144'hf11302d7fe7300f701a80a080137f912f69e;
mem[706] = 144'h0694ff04fefcfcb6f33af09ff628f874f883;
mem[707] = 144'hfe87066bff4d022e07faf41dfee9fca40d69;
mem[708] = 144'h0de7069a013cf87cf78a0dc9050ffcb7f305;
mem[709] = 144'h01c009f4fade05b803170dff086bf6620bb9;
mem[710] = 144'hfd4704d2f80df550fcc9f506fa80f3a9fdef;
mem[711] = 144'h01810b24f93aff22f40c015cf9a50e6ffb2d;
mem[712] = 144'hf28dffa5f308fa0a0c3f0f50fcc1f0da086e;
mem[713] = 144'h0175019b0242f25e0f530b61fa9cf60df253;
mem[714] = 144'h036607b6fa5bffa80f470698f5f6ff65f1d9;
mem[715] = 144'hf5630b26fa4ffa7c0ba8086704f0fbf70d81;
mem[716] = 144'hfac6fd41efd607bd01f9f32ef77a06a10847;
mem[717] = 144'h0f020ce500aa07090018efc204b4061bf8f8;
mem[718] = 144'h08fd07d00aabfe020146fa31f847fd71fb10;
mem[719] = 144'h0204f761fae6031af9fcf34efcd90ab00762;
mem[720] = 144'h0b18001e03a2fdcf0325fc8a04a00a61f4dd;
mem[721] = 144'hf4ddf9800dd401c7f3ab037cfaa4f25bf747;
mem[722] = 144'hfef1093301100c270937099bfb490e64f21c;
mem[723] = 144'hf254fb14f909f8acf6b305590f350903f0f9;
mem[724] = 144'h055fff320c0cff63fdb80ed5fdc800bb0e37;
mem[725] = 144'h05190116fc040ac4f62afa29f4d406010ae0;
mem[726] = 144'hfacffd480021fb6afe06fbc3efd6ffe2f5e6;
mem[727] = 144'hff4cf8440014fce50515f9b2f576f50cf7c5;
mem[728] = 144'h0bb9094bf47aff2b03350752f734f9c4f616;
mem[729] = 144'h0e2cf88e045e05f5fc2b0d500a31f072f23d;
mem[730] = 144'h01f7f975021cfbe00584f550037306f502ec;
mem[731] = 144'hff1905fefbef055c0969f380f967f795f675;
mem[732] = 144'hfe33fd8500e10c7b0246f928f7c6f09affd8;
mem[733] = 144'hfb59f24107440aaef3ab0b7e06cdfa19f441;
mem[734] = 144'hfaf60abffbd2f91509340c70f8c8f0fcf8ec;
mem[735] = 144'h0b3200bd0e200c2a09fd00a70060fe6a041f;
mem[736] = 144'hfb39fe42f4b8ff7f07b70235f5d90200efd3;
mem[737] = 144'h0d7a07dc08bb0e27f87af1ebfc1a02ccf938;
mem[738] = 144'h0b1e0ec7fe49078308c00b17070b0fdcf4b3;
mem[739] = 144'hf3b407c1fbc9f2520cb906fa0460075ff827;
mem[740] = 144'h0a84048307e703910926f43a06670326fd30;
mem[741] = 144'h0e65ff300eacff63f00bfa9d04290536f878;
mem[742] = 144'h0723063cf0f20ec1ff6804e8f298fc5b0c47;
mem[743] = 144'hf42101e9fc260559fde9f946f72402a60bda;
mem[744] = 144'hf337f055f36f0c5ef650faa3098d01400826;
mem[745] = 144'hf5db09690f560ccbfc2900950cfef967f96c;
mem[746] = 144'h0937f4f900160e060a16fcbdff6f0dbafab0;
mem[747] = 144'h02f8feebf41af857f83507090b820ed70ae1;
mem[748] = 144'h04f1f1c9fb06f9400e630db3ef8df67bfe3f;
mem[749] = 144'hff1806f105ecf7a30649efdcf5a10b20fecb;
mem[750] = 144'hfba50d50f46600c2f9850377fa7407c4fcf3;
mem[751] = 144'h049ffb0bfedaf433070007bbfb2cfe880bc0;
mem[752] = 144'hfd53fa95fc6f0bdc099208f5fc5403ea0aa1;
mem[753] = 144'hf2ca068a070cf7f2f51cf07af5dbfeff0ddc;
mem[754] = 144'h019903b4000cfaaaf086f261f13efbfc03d7;
mem[755] = 144'h0ac003ff0afaf264f0c906fb04010680faf7;
mem[756] = 144'h0860fb1d0cdc00a3efdf0cd009200ab2f7bd;
mem[757] = 144'hf8a50d880e2b097905b4f4f20dd900fb08f0;
mem[758] = 144'h06e80bd9f12700abf297f31df34402430137;
mem[759] = 144'hf173f65f07abffe0f3ee0ac3faf8055108b7;
mem[760] = 144'hfe17f2b9098305bc0755f2d0f7deefeaf7d3;
mem[761] = 144'hf7c20d2303fdf552f0720dcf04f30371fe70;
mem[762] = 144'h0f19f5a4fb9efb2e05310bafffacfce2f5b2;
mem[763] = 144'h0b260af5f793fa160d690c89f822f9e7075e;
mem[764] = 144'h0034f8b3093100ce05ebfe3ff6bafa26f4ea;
mem[765] = 144'h0a7b076202940b07f423fb0b0d5cfb0207eb;
mem[766] = 144'h08ceff8c023cffdc0b8d014907cd03dffce2;
mem[767] = 144'h0cfcf6caf91002bd0079fc76f7eef6960306;
mem[768] = 144'hfdc105340cddf8e7f328fb0bfbb5f142fce3;
mem[769] = 144'h0328f6730112007d04bc0188030df5ac03c7;
mem[770] = 144'hf7590d49087209caf7c50d4df051ff4d01ee;
mem[771] = 144'hfdf6f8caf7f8f1d20c270e52f49b0b5b0a93;
mem[772] = 144'hf2def357069508590a7cff0ff31dfa3cf7b6;
mem[773] = 144'h029bf55ef624f602fcd8fce8f8fdf446f04f;
mem[774] = 144'hf11e09fa049e096efa9009440406f47e0749;
mem[775] = 144'hf1cd01820e4a02e9f4bd015c0bfb016401f9;
mem[776] = 144'hf149fd0a025dfd9a0b73efc4fa5f070df981;
mem[777] = 144'h0e670b5df4b00f38f8d60fe1fcc3058c002d;
mem[778] = 144'hfdbcf0bdfd1103fe0fcd0eaef0690926fada;
mem[779] = 144'h0792086f05ff03b0f07209a10f29efcdf7bb;
mem[780] = 144'hf091ef9c06eafe0ef3700ccff1140b3a0bf8;
mem[781] = 144'hf3e0f475fe5b0124060f0763f1730ec6ff30;
mem[782] = 144'h0df1075cf823fa98f619fcf3f58402e70841;
mem[783] = 144'hf440029e0fd20e50fffa08a1f183fa47f3e4;
mem[784] = 144'hfc44045403aeffea0da0059002da0883fb13;
mem[785] = 144'h0b6bf07c01f60e59f9dd0efdf91f0702f7de;
mem[786] = 144'hf3dff40b053afaa9fb1709fbfeddfef9ffb9;
mem[787] = 144'h07840b0cfb490006f48efbe008bf09d0f048;
mem[788] = 144'h029ef7f8f8f8fc2bf5e7f69bf7d50c560587;
mem[789] = 144'hffb30f6403c1f3e9f116038406abf11efd6f;
mem[790] = 144'h02fe07f1ff3004d9092b067c03ba02d60e3d;
mem[791] = 144'hf9520f62f1b7f0b5f98ffea10cdcfeac0142;
mem[792] = 144'h01baf5c90c35034cf9b5f0ea0e70f29af86a;
mem[793] = 144'h0a7bfdcc0f56fd13f00e0aaff0d2f1db02c8;
mem[794] = 144'h0c8804ccf62af3440c2401fbf327f2ed02ba;
mem[795] = 144'hf88b08c7f1bcf215fa5af971f3750107f582;
mem[796] = 144'hf12cf577ff560c29fd43fad008260c33f20b;
mem[797] = 144'hf6760e780430ffbb0abcf19ff8440698f3bf;
mem[798] = 144'h0eb9f6b90574052bf248086cf60a032e0416;
mem[799] = 144'h0329fc1000b40d6df121f332fb2efebf0bb4;
mem[800] = 144'h0f350d940738f74003930a2bfaab0a5c0dc3;
mem[801] = 144'hf1e107a4f93cfd5df3ce0d9cf7550b27f217;
mem[802] = 144'h01b3f53af86ef662f2f6fc7af3aaf4bbf5bb;
mem[803] = 144'h02cc0cb504e5fccc0d9b0920f4d10a57fe7a;
mem[804] = 144'hfb34021dfe33f6db064af7cbfe830ea807b5;
mem[805] = 144'hfe780a9f0d37fba8f5e8080f05c30e14fb00;
mem[806] = 144'hf470091a04500d890b83fd74f4d4fee5fd5f;
mem[807] = 144'h05a207dc00f30a580339083dfa4a06dc0cba;
mem[808] = 144'hf5bc0a8df926fec3035ff07e0009f3c90b0c;
mem[809] = 144'h0874089ef332f91002a4050af6f6f19df1d5;
mem[810] = 144'hf2e4f7b70e7d02b4f3140623037df3b409c3;
mem[811] = 144'hffd6f0b9005af08c0986088ffbe2f960f945;
mem[812] = 144'h065601610c180a510b07f66e0ef2f571f066;
mem[813] = 144'hf7b9f680f910fac008b5f961f696fea50dc4;
mem[814] = 144'h0f0c0c960404037f0e2204e80aeefefafc7c;
mem[815] = 144'h0dc507adf77ffd650cedf7f3fcbb051b027d;
mem[816] = 144'hf445fd09ffa0fd17f852ff93ff0e0932f8aa;
mem[817] = 144'h0960fbfdf531f7710550f4e5f228fead0154;
mem[818] = 144'h0975074e0394003905effe6200740681fb12;
mem[819] = 144'hf512fe5b0e6dfce4f546f59bfec1f4760233;
mem[820] = 144'h0a8afffff5a60cb00e38f6550b44f7e50201;
mem[821] = 144'h08770358f230f7fef8e4042ef9caef94065a;
mem[822] = 144'h00740850f871f471f8ddff29f5cf00b20e61;
mem[823] = 144'hf6510e8b0d4b05bdfcd20a04fee101bf0e63;
mem[824] = 144'hf264fd420a2e076ef76e053008d606c30559;
mem[825] = 144'hfacf070ef812081e077ff2eefaf10a58f077;
mem[826] = 144'hf1e6fb54f192f877fcc204750716f4dc0374;
mem[827] = 144'hfc1cfdf90922fca0f290f6f2fc54060403fc;
mem[828] = 144'hfa22fb330dfef9ca046d04e70be8078bf4fa;
mem[829] = 144'h0183058df605fa58057509280bcdf58cf624;
mem[830] = 144'hf224f3b605a709a4f5b709200c81f3e60ce3;
mem[831] = 144'hf30a05b7fbbaf3cc0df30d9105fd0278f104;
mem[832] = 144'h01dcfad701e4058d024f00df0291f8480c7d;
mem[833] = 144'hfd1306be0cc50057f9fb070afa2804e8077b;
mem[834] = 144'hf526f6ee0fa10d0afb4e0ddb04b9fb23fefe;
mem[835] = 144'hf301f967f0880bd6015b08bdf711f33f0ded;
mem[836] = 144'hfe9909e7f3ebf41d06ec0f5defbef3fa0c30;
mem[837] = 144'h00bef4a1f427f2190280052a00ebfa500a4a;
mem[838] = 144'h0753f7d60661f162054ceefb019a08adf0b6;
mem[839] = 144'hf20f04d102a8f904f4f304fffb6c0cf10304;
mem[840] = 144'h08590bccfbb20249fce50816fa230a2af165;
mem[841] = 144'h0f1f0dc1020bfe5bf3d4ff1301bb078a0267;
mem[842] = 144'hf05efd9f0a59ff64f791f3dbfd5eff0cfb34;
mem[843] = 144'h0209fabcf267fecd01f800820613f0f20904;
mem[844] = 144'hf1c601b706e1ff04fbe1091eef57fd200553;
mem[845] = 144'hf8330c36f0d6f4670108f9ecf9f9f8da062e;
mem[846] = 144'h096e04900797f7b60984f809055cf3e804b2;
mem[847] = 144'hf0e60636f94cf3680dd8f51bf792f0860289;
mem[848] = 144'hf880f22e0e2b0060fc0efb8502f3f7f4fe5f;
mem[849] = 144'hfe7d0331f135f2050f1a01fc0548f7eaf1d5;
mem[850] = 144'hf57307f3047ff6fcf78b0bf9040b0465f279;
mem[851] = 144'hffc702dbf5a1fd4a0adff20e0b4d0cd9f3d1;
mem[852] = 144'h0cad06f0079cf688fe9df526064ffa9b02fd;
mem[853] = 144'hf8710224f06b076e05a1fa77022bf3e901d5;
mem[854] = 144'h0426f9bc0926f64202fb0be2f32af66c06e9;
mem[855] = 144'h0258052f0eba057cf38cf421050802d1042b;
mem[856] = 144'hf1590bbcfdb5f166043f01bdf1ce00eb0cf0;
mem[857] = 144'hf71c05a7f29e034eff4befdaf0a8f91b0e0a;
mem[858] = 144'h09df05fffb71f8bff173026ef37d0522f6ad;
mem[859] = 144'h069f01d3f61c042809d6044d0b500b8cf689;
mem[860] = 144'hf6310cfbf14909b0f082f962f766ef82f21e;
mem[861] = 144'hfae4012c0c3e0ee2f54ffe90fa6df0e109c2;
mem[862] = 144'h077700950fdd0527018e0aedf58906b5f646;
mem[863] = 144'hfa2dfe3bf9010b7b030dfbe50d340f3ff876;
mem[864] = 144'h0d38f787f09dfb95f225f67d094af65d09fc;
mem[865] = 144'h084509e8f101f1e00cb403b0f2000d5c0225;
mem[866] = 144'hf99cfbd1f57108bc004df411fc83f49af4b8;
mem[867] = 144'hf9b4fb45f85e0470ffc5fb34f87a02270d00;
mem[868] = 144'hefddf78c0077f5830f570398083f0f42042c;
mem[869] = 144'hf2d609df024ffd66f794f68603c6f0cafb8d;
mem[870] = 144'h0ee3ff6ff68afb550d7bfd91f808f7d30845;
mem[871] = 144'h0770041df46cffbcfff50dd2fbf2074203c7;
mem[872] = 144'h098cff5c062a0245fff7f4fc07d2f2710e49;
mem[873] = 144'h088bfb150b77f3f305c906b906690c77f11e;
mem[874] = 144'hf424fcdb085e073efba004b4f25af3e1f380;
mem[875] = 144'hffc6fa48f52df7a2f65201b8f31702bcfb25;
mem[876] = 144'hf3860dd9f46cf051faeefff1f582f2aff428;
mem[877] = 144'hf229fc91fe8d0d45f010ff7df1e00646fa48;
mem[878] = 144'h0ef7f691fe90fbd7f72403a706e20c46049a;
mem[879] = 144'hfdbe09c3001b00d9f13f0f95002bf182f664;
mem[880] = 144'hfd380890ff0cf06ef75501b402a4ff11f828;
mem[881] = 144'h031ff23cf65bf4fb0f1a0b56f74cfac4f5be;
mem[882] = 144'h067901a50a0809e5f83c044d0824f30d0162;
mem[883] = 144'hf8130139fbc308720c72017ef3e8f538f3ef;
mem[884] = 144'h04f6f3b10e36f991f3e8faf007c5f8a10429;
mem[885] = 144'h090e0bdd028005900d6afb6a063901b1fdfa;
mem[886] = 144'h00600eb3fb7e0027fd72f47df553f7aefc1b;
mem[887] = 144'hf7e00582058ef83b0d9d0348f3ad091bf674;
mem[888] = 144'h0e7801a0019005950692062cfd8ffeb70c16;
mem[889] = 144'hfec6f2320a1ffeccfb34f2b8ff20fd3df42f;
mem[890] = 144'h0bcb0e100542f7cff0730e53f1bff1360197;
mem[891] = 144'hf8650deaf88b001d02dcfc7a0100094c0539;
mem[892] = 144'hf2020b6907acfa69f0d6f4cefaad0a350acb;
mem[893] = 144'h06adef47f226fbbc084ff90b073ef8080310;
mem[894] = 144'h014afb7208eb03550025f725f7e00b90f359;
mem[895] = 144'hf1de0eccf6b9f6bdf1ee0ae500dc04d9f290;
mem[896] = 144'h0e070e72f46cfd730dc5f64501ce0452fd26;
mem[897] = 144'h0cf8f60907f50c0bf28708e4f0cf0b58fe94;
mem[898] = 144'hffe300830a10f2edf38a05380aaeff440b4f;
mem[899] = 144'h0a1bf0130663fdaaf34c00c3f107f1f8098d;
mem[900] = 144'h06800c2ff26e0f37fa59fea30e0af64af24c;
mem[901] = 144'hf7260b2effe20207f7cb087ff3fafd5fff50;
mem[902] = 144'hf63d0547eff20dc30b200fa7f6fc00940ef4;
mem[903] = 144'hfc47076904d907280302ff79f4d6f5d700ec;
mem[904] = 144'h064c0eb80ea409e201f1029ffc370c540c97;
mem[905] = 144'hf57d0d22f5300f65ffbcf7540e19ff15fff4;
mem[906] = 144'hf247f98d088c0a45fdc0f58305f0f705f1a2;
mem[907] = 144'hff1df4d3f2a609e5f0700ff50586f79001a0;
mem[908] = 144'hf87cf8ecf72a0dfb06eafd40f829f531ffc0;
mem[909] = 144'hf6a7f974fc9008930cb0f240fc80f3f903c0;
mem[910] = 144'h0662f65cfcdf00acf2cefe910829fb030ed2;
mem[911] = 144'hf831f3dff409fa96f77ff25300a5f25cf3af;
mem[912] = 144'hf2b8f05fffe9f0560df9f4a9f6f2f572fda0;
mem[913] = 144'hf70b0d710cf5069bf28bfd8c0e60f610ff7d;
mem[914] = 144'h06ce08720267000c07f503f3fbc00e3bf4ef;
mem[915] = 144'hf903f584f7ddf750f05cf1e9003df543095f;
mem[916] = 144'hfe23002d07bff4af0ef209a5faf906cd05e2;
mem[917] = 144'h0bc0f82efe0d0bd6f4c50463fc740731f735;
mem[918] = 144'h02a90e4f0a4f0a2dfe720bdd0d7904560ac9;
mem[919] = 144'hf7a30adb0734f1b5f189fd5505920abff972;
mem[920] = 144'h05cb0baef2f2f9100b740b93fc33014dfd40;
mem[921] = 144'hf804fb03fddb0fe4f2ccf8ae0e3c0770022d;
mem[922] = 144'hf2dbf5cc0804f4d5075c0858011ffa44070c;
mem[923] = 144'hf44bf3c3f77a0222033d04fdf8a3ff88046f;
mem[924] = 144'hffc900d3f54602c90478f26c074bfcf6feac;
mem[925] = 144'hf7aef965faf80c13fbc3f3c806e8fdde06a9;
mem[926] = 144'h0f4df9fc0483f3ef068cfceb0a40055100fb;
mem[927] = 144'hf23f0266fc80f7aff842079df168fa9d0277;
mem[928] = 144'hf25df2ad07b602e90ae4fddeff720ee80c05;
mem[929] = 144'hff85f9cd04ac0e950ef105ecfcd9f8d60130;
mem[930] = 144'hf134f39000160dfcff82fc65f178f40ff699;
mem[931] = 144'h0e62fd6bf8def1c7ffb00ce6f2470659f443;
mem[932] = 144'hf7800b90f5d8fc180bacfe1dfc04feaef865;
mem[933] = 144'h04fe0135f4570833ee7208b7fbff03fbf398;
mem[934] = 144'hf2eefa7f09aef658010ffbccf1effdf0f209;
mem[935] = 144'hf6980a090d8cfdfb02f8f6e4f590f50b0dc8;
mem[936] = 144'hf6af01b003d1095d084d0ac30a4ff0560b90;
mem[937] = 144'h05d20b720044063dfc21f8b301700bb1039f;
mem[938] = 144'h041e0885f1acfec90a4f0c4f0fa9f889f654;
mem[939] = 144'hf5bcf06e00f9f40d0f4002c6fded0b750f1b;
mem[940] = 144'hfc06fcdb08760460fb990d410545f0af09af;
mem[941] = 144'h0a5afccbfa91fafdf7380c4af610faa30bfb;
mem[942] = 144'hf4dc0c99eed0f2c5012cf6d60bd80dfdf46b;
mem[943] = 144'hf4e3f872028c077f0894023e06ddfc910d08;
mem[944] = 144'h05420fc5fa8a055a00c3062a01fb09830d5e;
mem[945] = 144'h065df80bfd63092b0031f924f61bffd0026d;
mem[946] = 144'hfc690f63fabcf3a2f1aafbc7f42305410d8a;
mem[947] = 144'hfbcdfa8f05a40f04078a0f2bf63df91a0353;
mem[948] = 144'h0cfc0f1b0beef21c0862fdca0a00fe930514;
mem[949] = 144'h0e070d4309f002560239f3fdf4d3f39df787;
mem[950] = 144'h087bff73f0c907bef1100e9f06640304f945;
mem[951] = 144'hf379f2260c6bf896feb6ff1a0b51f0adf15d;
mem[952] = 144'h0878f4e7f1d70e8dfadc0a32fe7eff0701c4;
mem[953] = 144'hfb44f311045b03d00335f677f646fe250aa3;
mem[954] = 144'h02400027f1fbf4760e10fae80c280d2ffd00;
mem[955] = 144'hf539f3d0f7ba015b0e8ff1f60fd3fbebff7f;
mem[956] = 144'h049d01d7f7a7f99709cefadbf18cf6f0febe;
mem[957] = 144'h0c660c61fe07f2f5f07bfbae036d047d0117;
mem[958] = 144'h0b44f655f68e04a70a870f6c0b0ef820f631;
mem[959] = 144'hf33e0b1409e909fa006303f00d91ffe6f8f9;
mem[960] = 144'hfa63f0600f1b04e40c77f3f1f0fbf86a0784;
mem[961] = 144'h02a607b101c7f1efff18f5a0f9c102baf392;
mem[962] = 144'h01fbfe1c01edf0ecffddf9c603730a32f844;
mem[963] = 144'hfaaa005defefffb6ff2c022f049af0d6fb99;
mem[964] = 144'hef95f82ff1a40bc7f1d607be04c9f2410e2e;
mem[965] = 144'h0468fa10f67b0b8ffe2af0af09c5f9a60cde;
mem[966] = 144'hf5390b2afb9800a800d9f66c0b29f7cb0ef3;
mem[967] = 144'h034cf358f914f86e05d4f8ef0b4b0b4a061f;
mem[968] = 144'hf3c6efb3fec60d1109e508cfffcfff7af2eb;
mem[969] = 144'hff4d0593f921070907f60a09060a08be0205;
mem[970] = 144'h040afabb073a0383f19d048f08b8f0b50070;
mem[971] = 144'h0ae8fffafd2ffd30f566099905fd0b27fc2f;
mem[972] = 144'h07d6f2e4f98007d30caa03f3fcb70eb4012f;
mem[973] = 144'h0d43f45706c4064ef8230f240ea30d8007fb;
mem[974] = 144'h0a43087ff82ffe5df9d9f1f00947f2dcf91e;
mem[975] = 144'h0beefa87fa4ff629fa07f000f3dc00e4fcbc;
mem[976] = 144'hfce3f52d0706ff26f1edfa47f7c6057e0e2a;
mem[977] = 144'hfbe1f2750f4d02e2fcfc0dc603daf0a5fb0c;
mem[978] = 144'h012bfdf7031f03d10090f3870adc0580f9e3;
mem[979] = 144'hfbbff7bff57ef21cfa9309a4f7bc06a5fc09;
mem[980] = 144'h0ce9f8cf06bb002b0697064bf54a05c0f921;
mem[981] = 144'h0d2af2d2f8b80d22f8f1f474fd6605ea0226;
mem[982] = 144'h0172f7abf72ffa770394f8d2f0fffc98f4c0;
mem[983] = 144'h08df040bfe67fb7c0dd30fa205f1f68b0251;
mem[984] = 144'hf8e40ba1f64df99cfd2cf9f0f21e0ae9f48e;
mem[985] = 144'h0cfcf16af20afc82fb9109dfff62febb0f43;
mem[986] = 144'hf00ff6470a2308c9fb27f3ca0a28f236f9ab;
mem[987] = 144'hfa6904590ebafcba05a7f153f6d5fa4a0026;
mem[988] = 144'h011700930f76fed4071c0300fff9f996058f;
mem[989] = 144'hf01100ebff6bfea9f9f5fafe04560150f83f;
mem[990] = 144'h0ea40d7af2a60555fd86fc59f411f16df8c7;
mem[991] = 144'hff15f3cd0b19f778f1010b040a5e0e35f926;
mem[992] = 144'hf300f0ed06f301910946ff4eff83fcb2f4bd;
mem[993] = 144'hfb17f4d4097a00ae0f92016109470f7bf30f;
mem[994] = 144'h0a6bf72dfc2e067c0871f97f04080b510d26;
mem[995] = 144'h01baf5b7046cfea9fa6ff89bf67008040f61;
mem[996] = 144'h0f9502f90bf702fcff8af745ff480dc2007d;
mem[997] = 144'hf14ef6f200aaf334fea20dfa0d7e01cff64c;
mem[998] = 144'h06cf055b0b03fbca06fe04db0d8c0dd3f18a;
mem[999] = 144'h052705ed00aafbc80e3a09210500f4d6f6de;
mem[1000] = 144'h0dcaefb5f180f073fc410aa40c48efe106fc;
mem[1001] = 144'h0fbf038607ff0ac30dc30bcf0c78f8acf20f;
mem[1002] = 144'h0f1801f7fd7605bdfa7ef99b082406ac042c;
mem[1003] = 144'hf574f0d504ce0e96f61f05d90683002505c8;
mem[1004] = 144'hfa12f259fa3703db0f70ffb7fc96fe78f55a;
mem[1005] = 144'h04caf8c50ac4f95cef720f8d0acafd64f0b3;
mem[1006] = 144'h0114007100cb012ef54bfe9a0bf9fe9b0dc9;
mem[1007] = 144'hf593f54f093b0d800f10064ef6840d880807;
mem[1008] = 144'h009ff3ed08a70349092d0930febe0f110d20;
mem[1009] = 144'h002e03760c9cf38f0da1ff9ff6380c9afd5f;
mem[1010] = 144'hfb54fa2008f1f9ac0708079bf41e0fdcf61a;
mem[1011] = 144'h009ffbc1083df3a00eb5f020fc2405a1f1bc;
mem[1012] = 144'hf0b403d4fd07f78c00870cd5fba70c9b0b88;
mem[1013] = 144'h0d11fa93f856f14108fafbea068307bf0a40;
mem[1014] = 144'hfb6af0c20cd2fdce017ff811fab5f2bcff83;
mem[1015] = 144'hf954eea0f0f5f90b00c703a8021ffb970e7f;
mem[1016] = 144'hf089fb0bf9c6f2f1f97c05340e2f059e0b79;
mem[1017] = 144'h0c810c380fb2efee0d45f2370ced0fb2071b;
mem[1018] = 144'h0c1c08c5f2a6f8a1f584f339feb80326fe6d;
mem[1019] = 144'h0d25fa340e3ef1e5f810fb89f32c070908cf;
mem[1020] = 144'h074b05dc0d1bff2f03870790f2b1f5670043;
mem[1021] = 144'h0be706da0b9af0bf06aa039308140088f00a;
mem[1022] = 144'hef92043ffa94f39efa85f9b20b77f9f50dcb;
mem[1023] = 144'hf463fb8b0ae00beff800fb72faa109b203fc;
mem[1024] = 144'h0dd4ff6afdeb057cf5aef4f008a7026df801;
mem[1025] = 144'h02b9083b0e050df8fe0efc75f6f4f3170c15;
mem[1026] = 144'h0975f72e0f89f30b0752f398f225f8db0087;
mem[1027] = 144'hff91073f088604670c530f33f9f5fadc0dd5;
mem[1028] = 144'hf9ecf880fcf302f4f5c40030fc2001d70bf7;
mem[1029] = 144'h09d20e54f94d05c201e700def0f7efe40de1;
mem[1030] = 144'h0c8ffc600acef5d2f2a8054df671023ff13b;
mem[1031] = 144'h002afa8cf391080bf056f77403d3fd37fdbc;
mem[1032] = 144'hfe2bf5e207bc04b2069703b1f824fa9b0615;
mem[1033] = 144'hf708f0c80280fce3fb22fcf503430afd085f;
mem[1034] = 144'hfc4309cc0c2d0352f365f56e009f075a0455;
mem[1035] = 144'hf7a5f79afeca04800a5601c1f1b80cef0861;
mem[1036] = 144'h096dfa1c0ebf0647f4ddf5830196f2f608fc;
mem[1037] = 144'hf1c7f47b0ec9fb76fad90c8c0c0c06ce0e47;
mem[1038] = 144'h00aa0c9a0181fe0f0142f36b01370c1f03c5;
mem[1039] = 144'h08290f2e047af5f9fdbc0a7a01a9f102f358;
mem[1040] = 144'hf6a909530dab038803c6f051082c0cb6f124;
mem[1041] = 144'hf3befdf0f2070a41fc2d02fd09e5f17cf7a9;
mem[1042] = 144'hf9070dc500cc03790624f2c90e12f283fb6b;
mem[1043] = 144'hf7570f36075f0123fa9cf68d0285043d0085;
mem[1044] = 144'h07e6fcf6027f005e0bbbf49cf1720caafcc3;
mem[1045] = 144'h02c8f51ff3a70b38fde4027008d5f60cf963;
mem[1046] = 144'h065dffaef1fa014b097af55efd03fb8cf5ff;
mem[1047] = 144'h0b100ee5025800100274072704f8060ef9db;
mem[1048] = 144'h0cc7f04505b00d190cadfc7b0eaa05b60486;
mem[1049] = 144'hfa83f5660f75040b0872fbeef4b10041f944;
mem[1050] = 144'hf86ff0c70dc70ed70bac00a9f664f014fdce;
mem[1051] = 144'hf586f8460577f263fb72fb56038ff37402e5;
mem[1052] = 144'hff05fa5b006f03c70c2903d6006000b1f6a2;
mem[1053] = 144'hfd73feb6f9360945fe900041f040f86b03a8;
mem[1054] = 144'h04f7fbddfb93f46506d9f530f1eb0bb7f35a;
mem[1055] = 144'hf3b8fcfbffd805cf0b3c015d0c4ff5bbf39a;
mem[1056] = 144'hf2b9f52902c6f4dc06430d2cf0c2f71f0c2e;
mem[1057] = 144'hf86704f7fc24fec30de9f201f8950eb2f72e;
mem[1058] = 144'h0f89f00bf077f3d8ff60f9da08bc05f0f35e;
mem[1059] = 144'hf11a0818f7dcf1fffd39f2c0fc54fb6ef697;
mem[1060] = 144'h0f58fe130023f7d3f8b1fff3f6d6f259f981;
mem[1061] = 144'hfdbffaf1f6d30af30d8bf030f2caf973084f;
mem[1062] = 144'h086d0a7702dcf2fe0765f58bf18600190bdb;
mem[1063] = 144'h067707ca031907ed04ac0cd2f5fcf710fa8b;
mem[1064] = 144'hfe26f2abf7f60b8efce3fb7d00b3fcc6077e;
mem[1065] = 144'hf4d6fa260445f49ff1b2ffd9029ef687f594;
mem[1066] = 144'h0417f759fd63f8b10ad500550863019707c1;
mem[1067] = 144'h0c760bc702b5f5c1061ffacd0e8ef86403ec;
mem[1068] = 144'hfca804920accf844f1f0f9a905cefb4a0289;
mem[1069] = 144'h008ff7d109cff39c046f0e71f88dfbb9ff8c;
mem[1070] = 144'hf1b1f8f9f258f9b5ff090043f8320abb00df;
mem[1071] = 144'hf5570dfe08f70d4df6ae00cbfe1b05a6f89a;
mem[1072] = 144'h0d200686fd0ff7fd05cffcbf021defe5fcbc;
mem[1073] = 144'h0388f1ba0d4703a104fa086706b8f75cfe0b;
mem[1074] = 144'hf8d3f2070296091e03edf9ce00acf1a503d8;
mem[1075] = 144'hfe2cf4910668f0ebf47004f906cc055702ee;
mem[1076] = 144'h00adfdb0092903da0d160eb7099304b40199;
mem[1077] = 144'h01b2f45604c8083904470897fbdf04c10bc9;
mem[1078] = 144'h0aff09db06fff6e805fa0885fd1e07b0fe48;
mem[1079] = 144'hf4a3f7f4f09f03c0effd0036f9650dd6061f;
mem[1080] = 144'hfc31f56d075efbda0576fc90fa1d006602bc;
mem[1081] = 144'h07200a95f92cf72ff3850d0f05d003180f1c;
mem[1082] = 144'hf40d098afa12fd540a3a02f7f5d403dcf7c8;
mem[1083] = 144'hf70df4700f81f012fc1cf12efbbcf64900f8;
mem[1084] = 144'h0106ff680e060600f546062e0e7df0560f48;
mem[1085] = 144'hf674ff45f7ae09a40193f3fefa1d0777ef5c;
mem[1086] = 144'h03b0f509f1f204240241f4db0aec0d8e0312;
mem[1087] = 144'h050304320161fe06fb28ff73fbba05410532;
mem[1088] = 144'hfcff03b30644f1ab01adf8af02d00dac01a2;
mem[1089] = 144'h087c09bc0b8af44a05270822f3b9f86604af;
mem[1090] = 144'hfb8f037af428fcfaf3340a520e3df4630b0c;
mem[1091] = 144'hfaebf58d03350a880d3a06a600d207e3fc8f;
mem[1092] = 144'hfac0fc090a83f468f9730f5906d0f598fa4d;
mem[1093] = 144'hf1b2f26302e3fc19f7ccf322fe6e083ff12b;
mem[1094] = 144'h0855f61b081f08caf362ffb606a90227f484;
mem[1095] = 144'hfe1cfc4ff605ff04f7f4f1520ccf09dc039d;
mem[1096] = 144'hf412f3c90308f41bfb5afab4034a03e4083d;
mem[1097] = 144'hf996f28bfe09f9e608d50a59fa72061df1b8;
mem[1098] = 144'hf7ec0c79f94400a6fa4af464fde0058df1fa;
mem[1099] = 144'h0ef5f418032a0433fa6101b1fbbeff3ff725;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule