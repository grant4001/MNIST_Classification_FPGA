`timescale 1ns/1ns

module wt_mem4 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h040f069ff0a702c9fd6df7b1f6a20dc4ef0b;
mem[1] = 144'hf47e0511f06ffaa8f7320db60312faa6fd5f;
mem[2] = 144'h073b054df365f370f9b8003f0ce5f286fcfc;
mem[3] = 144'h0aaafe0105770517f9cd03f20d2c08a00cd1;
mem[4] = 144'hfad2f79e09e8000d009102ec02b3fc3bfdd1;
mem[5] = 144'hf7e500d8f23004be0e4a0ab50836fb23f15d;
mem[6] = 144'hf39108c70723fbd6f60ff10efc53fc1efd8a;
mem[7] = 144'h06e90d38021bf397037e078c0511f1d2f60e;
mem[8] = 144'hf4e4f72004e900540ef7fdb20c220e19f523;
mem[9] = 144'hf4a1f9b7f2abf5c30b61f286f8af0529f881;
mem[10] = 144'hf1e6f3e2f94cfc8bf73408d6f5bef6a0029e;
mem[11] = 144'hf6470abdfae10497f6b2f0de0ac4f2a3f724;
mem[12] = 144'hf22803d0038f0815f3510acf0784ef950dd6;
mem[13] = 144'hf09c07ed0bdaf2f20513f0c306a1efe0081a;
mem[14] = 144'hf8910ec6f8180ab10055f367f022fb4d01d8;
mem[15] = 144'h092e0adbf49001e3ff33fdf6f24cfe41f527;
mem[16] = 144'hface0cb90acd0a9d009af81609ef0921f066;
mem[17] = 144'hef98065cf233ef410ad6fe3b0f490535f036;
mem[18] = 144'hf9a7ef51f2f9fdc2f967ff88fc2cf487f5ad;
mem[19] = 144'hf903f7e1f946f400f73c03a4f5fef66cfc41;
mem[20] = 144'hf46afd42fb6e0ac9031e099afd69040d0b7d;
mem[21] = 144'hfed0eefbf1c4f6c30279f44cf78e09ddf5ce;
mem[22] = 144'hfea50c1c02d2f261ef6c07cffc69f8cf0c66;
mem[23] = 144'h0bb6ff60fe9500f5011d0eaaf5c4f333f419;
mem[24] = 144'h0001fd260b3e02030e47fb5bf5000d76f16c;
mem[25] = 144'hf8bff7ca01620955f87cf6e6f0dbf1da06a5;
mem[26] = 144'hfe67f8e801810b39fc8107df04880c9b095a;
mem[27] = 144'hf21104c4f29def62f395f3060c54fd6efa44;
mem[28] = 144'hf63afe3f0acd00c808bf0aeb00a5fe26f1e6;
mem[29] = 144'hf251f8260e5a067afe86fed00b1707e70217;
mem[30] = 144'hf21902930863f2f0f9fbf29304b9fd2efc6e;
mem[31] = 144'hf26207e00ca90381f74f07d4fea30eac0969;
mem[32] = 144'hf6e1f731049effedf1adf6ed06cef97f00fe;
mem[33] = 144'hf6a7ff94f96105fafc060103f5eef3270920;
mem[34] = 144'hf5970ec6066cf13af6ceef7f059ff8f20c70;
mem[35] = 144'h0cc0f69b0b5bfb0508b205450130fae7f812;
mem[36] = 144'hf563ef5909ddff9d0799ff1ff3e00823f335;
mem[37] = 144'hef860a2fff890015fe840b820dcffbbb07b6;
mem[38] = 144'h00450acff35d0d4d02ef0db7080201ca0efa;
mem[39] = 144'h0a070dbaf1f0f32403680eb0073e087af0b8;
mem[40] = 144'hfef9f9b6fca2f6fffac8003a052d0423f38f;
mem[41] = 144'hfac4f8c2f95cefff0d39f462f8e202820c5f;
mem[42] = 144'h02d208d0ef3c0116f0870e2903a30a4bf227;
mem[43] = 144'hf1cef0db00530144f0f5fe15fe2cf802f637;
mem[44] = 144'hff280c40ef740cebf3ba06960bf20c5f016c;
mem[45] = 144'hf403efb6f2befc16fcb0fdb2f60ff71d0e12;
mem[46] = 144'h04bc0120f7b1f7870059fbe80e9707a50566;
mem[47] = 144'h02380a19027b0219f5c2fc910294ff5707de;
mem[48] = 144'hf76508f50dfafeb70beb0c6605da034d07ab;
mem[49] = 144'h00860ee1f1d9fc6a05840140f2f1fadbf98b;
mem[50] = 144'h046d0954054e059102eef7000a3403220537;
mem[51] = 144'h06ac0e03efdb0bd60833f00c0ce1f28f0097;
mem[52] = 144'hf9b9f94409a20c83038808ccf589f4cc0ace;
mem[53] = 144'hf07c0ec30bb8efa201d2089308e1f2040d22;
mem[54] = 144'h0f44f71a0b38f2b9024b00000edbf8950e98;
mem[55] = 144'h07c7f5f500dbf9f0f33cf3230004fb550e2f;
mem[56] = 144'hfa15f908fb1e056df163fe5f05d5f784f41b;
mem[57] = 144'h01e5f5df05faefd50594f83df361f2bfef36;
mem[58] = 144'h00870b92f74d099b0458efa203fd016e05ce;
mem[59] = 144'h09f8f206065f0bee09d9f87bf2d9059cf607;
mem[60] = 144'hf9db0158f09fffc80b29faa6efcdfb1e08b9;
mem[61] = 144'h0213f50b09eefbadf48c005f0c42f8d4f294;
mem[62] = 144'hfc7e053af27dfc2b0671093604ee08c70480;
mem[63] = 144'hf918fd48f3e3f0e4f813fe7b0739f5140804;
mem[64] = 144'h02b900ecf7bafa650bacfa43086b0259fd45;
mem[65] = 144'hf009f7e0f0dafdb6f50ef64405ca0a2709ff;
mem[66] = 144'hfe9a0eadef91fed3f05b0c000e5807a5fda1;
mem[67] = 144'hff6ffce905fef96efed3031a06fefe820e39;
mem[68] = 144'hf6550a0fff44f64cf581f9c30dfbfbbef8e8;
mem[69] = 144'h06a30af60e3302bdf2270a4e035df900f8c8;
mem[70] = 144'h0e63f1d8fc5e0df900e80543f9ef009efa22;
mem[71] = 144'h0b46f49ef5420311fb74fc73f3fbf93cefe1;
mem[72] = 144'h0c27fd32f8d90dfa0f5b0a890dbc0168ffc5;
mem[73] = 144'hf9f404ebf1a1f34bf6a40a47f16e0d8206a6;
mem[74] = 144'hf63b0e6af897f0fc0563086f0d01fdbe0e0e;
mem[75] = 144'h0557041403acf52f09ecf685006108ac0e33;
mem[76] = 144'h0cbf0d16027cfbc7fa56f6bbf85b04b40e0b;
mem[77] = 144'hf2290c41f0f20e57020ef14ffe38f5cc032b;
mem[78] = 144'h06b4023f0e36f50909b002f1fccf06a60e88;
mem[79] = 144'h0c130cde0a6f0c430c8af2f3fe9d00730db2;
mem[80] = 144'h0f760782f3a8f78afc710ac6f2070f2bf1a0;
mem[81] = 144'hfa8c087900530016095c0140fed00c2a0b86;
mem[82] = 144'h03ba06f9f74501f9f098fc21f0890667fdba;
mem[83] = 144'hffc8fbaa0979f85ef70f082df93ef6d705a5;
mem[84] = 144'hf1970cd6090cf4bd0ec7fa4b045ffdc1f265;
mem[85] = 144'h0e340140f56e0e810e4a032209800f4b0c93;
mem[86] = 144'hf71cf724045307760830f7c6f79a0156f34f;
mem[87] = 144'h00c1f698032b0e270928f839f8bef5bf056e;
mem[88] = 144'hfe05f0b80d840748f2ba02a2f79204ed0b8a;
mem[89] = 144'hf1e5f3a6effe0c4dffdef3010ac5f88d015e;
mem[90] = 144'hfb6af12c00a60e6dfe9f0b37f4f50340fb75;
mem[91] = 144'hefb9fb61fdd5fb7efa32fc580cc7f543f36f;
mem[92] = 144'h0375f52200530d2b00fbefb3fd03f3a5f5b8;
mem[93] = 144'hf4900d83f9a602fa01dafef4f2140c520c7a;
mem[94] = 144'h056004a707cff770fb9b016bfdaaff4b0c4a;
mem[95] = 144'hf8650f6004e80a37fda10e70f0540237f42f;
mem[96] = 144'hf2e30a88f02df433f9e1f9a9f8150037f547;
mem[97] = 144'hf996005f079d027707400c550710f5b7f34f;
mem[98] = 144'h0f44fdf30671f737030605f10f420694f7ec;
mem[99] = 144'hf843f213f13efed0f2de064f0e730260fe80;
mem[100] = 144'h03bbfe2f02d2f18e02def1affce4fa30f869;
mem[101] = 144'hfdfdf50c0e300d4bf70806f10fa5fe170066;
mem[102] = 144'hf714f694fafdf93a0afdfe5f077f05ddf452;
mem[103] = 144'h027907e80e0ef22ff0b6fbee099c0003f116;
mem[104] = 144'hf351f647fa4ff8d00280f0dff51a08dbff65;
mem[105] = 144'h0bb2f1c20d32fb1d0f9f080207d6059c07e5;
mem[106] = 144'h0f94f646fe3dfbb70a8af0c6f1f2f7a8013c;
mem[107] = 144'h0b9bf9f3059aff6ff7c9f323efac042bf8a0;
mem[108] = 144'h06500484eff80185fae40a480606f59a0402;
mem[109] = 144'hfa63f9f601420d9bfaba0d9ef6d007f3fb8a;
mem[110] = 144'h0e870e4e0855f792f53df299f3aef211f82c;
mem[111] = 144'hf4aa0900f6bd0d2e0b460052f621f1c604e0;
mem[112] = 144'hf14bf255f5ddf9e7068206f5f7f707930c76;
mem[113] = 144'hf071fcc80768f06af7d70c17f4c50c450794;
mem[114] = 144'h0cb3f859030b0eb0fd87f07a01c7fd8f01b7;
mem[115] = 144'hf37208310b60fcfb0bb4f02d0ab50f81ffc2;
mem[116] = 144'h070f0dfe0c6c061905b6f269ff9cf0fefb0a;
mem[117] = 144'hf9cef404051efe0bf83c004b0b8a0d6ffe2a;
mem[118] = 144'hf2b1062dfaed01b1fc8aff0701d500b0f89c;
mem[119] = 144'hf3cffae00ae0fedff41ffeb60dd10b150a38;
mem[120] = 144'h06db0cc7f04e046b003d04e006220a9ef912;
mem[121] = 144'h0deb0011f93ff13e004cf654f88509c3f1f9;
mem[122] = 144'h093ef561f849f8200c41012f08f0efe7fd39;
mem[123] = 144'h0e6b0a930f0c025c0e9efe380f31fbe6fbb8;
mem[124] = 144'hf0c5fd3e05f2faf3023df3acfb820620fb9c;
mem[125] = 144'hf467efbe0a3b083e001d099a0207f12cf2fe;
mem[126] = 144'hf3430485fe14f2d1f535f207f2c500cbf81d;
mem[127] = 144'hfa43f89df53b0863fe4ff8e0f78d0e4c0ceb;
mem[128] = 144'h0a8204fb0469f93306b5f2fcffec03aa0d3f;
mem[129] = 144'hf50e09b3078cf458087405fafdf10f45f96a;
mem[130] = 144'h0543fc250c0df7d80cc70327f2eff49d0c3d;
mem[131] = 144'hf03c095403560483026cf1d40d65f0380169;
mem[132] = 144'h0ce3fddef16e07b10e330d6a0e5ff26e09a5;
mem[133] = 144'h05180880fe63f5f1f8e0fdebf374f0be0c83;
mem[134] = 144'h02f90dfdfcdff8f90cbd0d01fccbf093f5b8;
mem[135] = 144'hf72af30ef861f6560cae01ef0201f21108e7;
mem[136] = 144'hf3ff0f0a06d2f028f8c7f524fa4dfd8cf9e2;
mem[137] = 144'h0f2a0ad30fc9f39f086a0b90f6ccf1d9f537;
mem[138] = 144'hfa2f039ffe5d0f2ef59cfbbd030ef532088d;
mem[139] = 144'hf7e6019303e7f3f1f789fc49f2da06d80fc6;
mem[140] = 144'h0e91fbde0bb5fe8102c1fc4706e9058b04ee;
mem[141] = 144'hf9e7fd8df4910988fb280d74ffdef9bff2f6;
mem[142] = 144'h0e19f9f4f584fc3cfbfcf2a508390ad7015e;
mem[143] = 144'h00ad05f60ae70dbdf8480b8903b5098b0599;
mem[144] = 144'h0c210cf70c150002fa38fc2a00a00343f29d;
mem[145] = 144'h0aff099d0d43f51c07d903fdf77905e4f0e3;
mem[146] = 144'h089b000ffded086304dff9bdf2460f49f979;
mem[147] = 144'hf7a7f4fe0151f77a0253f016069e08a6f367;
mem[148] = 144'hf598fcdc0ee905f20101f5030e4c0a7cfa74;
mem[149] = 144'h00d20b5bf835fe530d96f6200817fa56fa4b;
mem[150] = 144'h0280f6c6fc09013afdd204e6fbc8ff92fada;
mem[151] = 144'h0747fdc2f161fcbaf821070d02e7f0c6f548;
mem[152] = 144'hfb08005908b3024a08230cf1034e0363f4a4;
mem[153] = 144'h0a6906530bda010e08c3f9140e99efcbfb8d;
mem[154] = 144'h04f501a60c4af9e50131f51bfad40140074e;
mem[155] = 144'hfb74f2a1f80d0a2dfa4afc350b8a0b31f151;
mem[156] = 144'hfcf900dd0ac50ee6f63c0072f10f0c790f5b;
mem[157] = 144'hfa1e00840dcc0f98ff5a0a1308550d19034b;
mem[158] = 144'hf606fd9ffc67056cfcdff0b5fbf2fee3f8f1;
mem[159] = 144'h099ff075f917f16c0cafffd20ab8f39104b5;
mem[160] = 144'hf6bc00e4070d096208ed04040d88f887f119;
mem[161] = 144'h00df0207fa84fe9f0d7ffc42fd02f11f0168;
mem[162] = 144'hf300f8aa046f011f07660699ffbb0d3ef166;
mem[163] = 144'h0fbb01b6052df7580f300164ff0304b6fc6a;
mem[164] = 144'hf27eff9efa480060ffb7f6a10ec7f2adf1d4;
mem[165] = 144'h00e1f47df7520f51fcb00e3bf67904c30f17;
mem[166] = 144'h09b102f50dcc05fdf3a3f3ecf3bf0052fb0d;
mem[167] = 144'h0f930332034902bbf3c10def05b7fc76002d;
mem[168] = 144'h09c90b6205f107a0ff56f0f0074204fdf829;
mem[169] = 144'h0beb0803fbb1f1ac057402ebffcb0605f822;
mem[170] = 144'hf07708b401d9f47cf97dfbaa00cff6cc08d0;
mem[171] = 144'h02dc03ba0a3605ecf7d8f1adfbf8016ef7f5;
mem[172] = 144'hf8c2f665f6710e50f845f8eb026508b6f1fe;
mem[173] = 144'hf22408f7f7c706b1f037fa180896f15a013d;
mem[174] = 144'h0f71f9b40f1fefde07640d6af4640681fa54;
mem[175] = 144'hfa4f083a0c9cfe26f053feb70a06fc390f0f;
mem[176] = 144'h0ee1078c0aa6f02b01e7046efd15f390f357;
mem[177] = 144'h0132f0f1f772f598fe1d00500233f9eefcde;
mem[178] = 144'h043ff9a8f9a109a20b65fa2e0cb608b60e8c;
mem[179] = 144'hfc0cf7f2fceeff10f9c806defc54f6f7f37f;
mem[180] = 144'h0dc0096b00e6043aff74ffbc0efafae8061e;
mem[181] = 144'h0e76f599f528fa610e31f50afa9afff80add;
mem[182] = 144'h08eb0dedf18b0220057503cef999f4f5ffce;
mem[183] = 144'hfdeef154f4bf0ec70b9c0383f037f51e0042;
mem[184] = 144'hf492023bf7e4f074f0460ce3f8aff0d8f108;
mem[185] = 144'hf3b5f947f324f1b30c90ff83f6a60274fd29;
mem[186] = 144'hf9ba0271fb34025b0c870291fab5fadb0d44;
mem[187] = 144'hfb9defe8025f0ea4041cfa90089c064f03f6;
mem[188] = 144'h0e07086207dbf21cf8110e0500020bf8fae5;
mem[189] = 144'h0c1cf00b002c0653f508f0d809a2f8ad0108;
mem[190] = 144'h02a6f1b4074b099c02530fc80436f553ff86;
mem[191] = 144'h0586f0ef0a980e9efc16057ef761f4e50d9a;
mem[192] = 144'h0afe0462fb4d0b8bfe4c0bf2f47c01d0fe37;
mem[193] = 144'hfc5f0c92f603f654f760f0e8ff10f9b000e7;
mem[194] = 144'hf5f7fde0f562ff8e0eecf6f005f60356f717;
mem[195] = 144'h031ff3c2079e0ebef4600eb0ffd40fabf47f;
mem[196] = 144'h0903fc53f10c0805f313034f0a02f02e0b9e;
mem[197] = 144'h00f2f53d00e4f63004ddf7fa05e705a3f196;
mem[198] = 144'hf145fa46fb4cfdc90addf26e03f1f2a8fa2a;
mem[199] = 144'h0743f5c5f1f2f85a031e07e2f3d5f9840797;
mem[200] = 144'h077305cc023e091df4a9f9450d0a01270d86;
mem[201] = 144'h00e0f3a0fa4c0a00f06a026c08c9f75c0e6e;
mem[202] = 144'hfd0ef0e9f39502b0fd550a64f63bf18ff9ba;
mem[203] = 144'hfd2a08b60502f0fe0d95fb400cfbfc3508d1;
mem[204] = 144'h04bffa23f84602d4fd8c0569f4fef70d04ac;
mem[205] = 144'hf196f36ffb0efb5a0ad40fae0dca0080f744;
mem[206] = 144'hfe6403470ae7ff790c8ff284f88a0a680a67;
mem[207] = 144'hf978f3cbf4d909740288035c062f072bf9d7;
mem[208] = 144'h085cfa040f280c81f31df1cd04fa0e4af404;
mem[209] = 144'hf12a0642f8a8fe07021ff11bf245f6edf436;
mem[210] = 144'hfadf05fd05b9f909efc9f4c705b4f95b064a;
mem[211] = 144'hf5cbfa65f8570887f57c0bb40e7ff707f716;
mem[212] = 144'h0750091105d9f239068403c3f6e4f780fb3b;
mem[213] = 144'h0aa0ff0509e1f24bfacf076cf172f8f7f6a4;
mem[214] = 144'hf5d70970f8090c6bf8910e4f03be0c3f0156;
mem[215] = 144'h03ad0b87095b079c0a7e0cbe0e93f69bf5a1;
mem[216] = 144'h0ab701a20e4d0cfe04ee02e6fb84f9def98a;
mem[217] = 144'h0f97f96d0a410a9a071dfa7303e2f18e08fb;
mem[218] = 144'hfdeef34bf193026affb104030d5703ad01cc;
mem[219] = 144'hf122f968f9f9f4b8f2cd08f7052c0bec0aa0;
mem[220] = 144'hf31d0676007ff42a0b50f720ffbe09a0fedf;
mem[221] = 144'h0e4502380432f446fb67071d0d22f5f3fb2a;
mem[222] = 144'hfaa5f81ef1bbf2200c5504fdfa2ef2740876;
mem[223] = 144'hfc8afc7002f7ffbf0f55efb70dee03fdf5cc;
mem[224] = 144'h037902220b67fdaffd76f4810ddd0de70a6a;
mem[225] = 144'hf2befa52f27f096efb0f0178ff6bff6906fd;
mem[226] = 144'hf9d60532fe980007052702d2f9ecf01bf1de;
mem[227] = 144'h0f9ffbdaf51a027bf6aef865f651f92d0883;
mem[228] = 144'h0301f323ffcbfbd3f0bcfe68fdad0af7f85e;
mem[229] = 144'hfe4e0fd108390183fa9cfb2f08f80a9a0c39;
mem[230] = 144'h0576fbc3f4d004f602aa0a78f5bbf088042a;
mem[231] = 144'h017d088001f200e2f8bd067d0df1f8340b9b;
mem[232] = 144'h06c0fa07ffdc01edf437f1a0f1ba09c1fccd;
mem[233] = 144'hf98a0e680cdf023306ef066c07e7f196f1c4;
mem[234] = 144'heff3f24a031ef015f534fff3f9550ca904c3;
mem[235] = 144'h0e3dfb87f9040458f59c063b027d06f3f420;
mem[236] = 144'h07190c36073ff5d7fc3c0310fd9c00c4fff0;
mem[237] = 144'hf57d033ef7db0419fb300906fa04fa47002a;
mem[238] = 144'h03b4020c048bf5f1eff7087bffe8f79807a9;
mem[239] = 144'hf736fc13ef77fd0afd5c06fe0d490cd8f7ac;
mem[240] = 144'hf00cf2c50a63fa9efc9ff467f351089c0bd7;
mem[241] = 144'h06c20ea3f3f7f713f0070129ff9af7ac0c86;
mem[242] = 144'hf35afb2dfd79f41e0dc80805f22ef42200f2;
mem[243] = 144'hf0c301920682f632020bff9d09e5f1020899;
mem[244] = 144'hffe80869090cf2f80a74f022f438f5f703c7;
mem[245] = 144'hf6aaf7fef8740ee90e13f3a7ff9706860afc;
mem[246] = 144'hf56cf817fe020c20048b0a94f84ff5e00813;
mem[247] = 144'h0e8f03a9fee706e909d20f60019a0dbff13f;
mem[248] = 144'hf29cfbcb0cf9ffa9fbecf4b00650f8010f00;
mem[249] = 144'h0bb0f86d095806d0fa67f2f7fd36fa06fc1e;
mem[250] = 144'hfb5af41ef5b10617057e0978fa410815f8da;
mem[251] = 144'hf8edf9fdf272fd410dccf6a0f8790b13fe48;
mem[252] = 144'h00520ad608c2f2fff106f23e02c8f306fb92;
mem[253] = 144'h05fcf01ffc660251f7cd01adf60cf921f911;
mem[254] = 144'hfa93f71ef75707a6f7640bb8fa2a0565f940;
mem[255] = 144'h0dd90d1a0d06f4dc09f2f7ddf151f7b30efe;
mem[256] = 144'h0e0f002d0eb009fd024d0682fb2bf28e0f5e;
mem[257] = 144'h040f07eef243f0aa09def4b30ceafa550133;
mem[258] = 144'h0e400152f7a1f932087507dc0c0b0de6f984;
mem[259] = 144'h0c3afbedf5c003daf15ffd12f6cbfa9e0144;
mem[260] = 144'hf9f3f648040af28bf3f3fc7606a2f3de09d7;
mem[261] = 144'hfe2d0739fb5201c9f865014efc83f4e90e37;
mem[262] = 144'h00e40744f2fe000d0f51f571fe4d011707a7;
mem[263] = 144'hfe0e0bbafbabf89104de04d8efbaf61bf4be;
mem[264] = 144'hfb25f9c8055ff4d8ff53039603d6f9f8f851;
mem[265] = 144'hf65f0f8706fd0a33057bf70207f5f8a50a8b;
mem[266] = 144'h0b6702cbf141f9ebfcfc0dae0a4507d4f604;
mem[267] = 144'h08c7f6c90828fe83f3d3f11a0879ff3bf36d;
mem[268] = 144'hf74cfe29f9330599064a07def27503040924;
mem[269] = 144'h06ff08f1f98efb4f0574f1f7f3fe07080eaa;
mem[270] = 144'hf6c7f2ce064ff240f01d06a6f867f588f71a;
mem[271] = 144'hf64604d4099b094ef281f14af25805f7f7b9;
mem[272] = 144'h0269f3efff820dc0f2d8f054fb49fd9afc14;
mem[273] = 144'hfad208a70f91f7ad0d55029ffdce0f0c0361;
mem[274] = 144'h0eeb0538ff00041bff30f41b003df937f93d;
mem[275] = 144'h0da9f23e03310000f00d0d310d66f5020e0b;
mem[276] = 144'h0ddc0f7a03edf6d60d5b008a083e02af0de7;
mem[277] = 144'hf99d0395f99dfdce08f2fe7ef099fbf00468;
mem[278] = 144'h00660a52f178ffbb0f8defddeffbf0a00ac6;
mem[279] = 144'h02660ecff810081af7600ab4f2aafadef7cd;
mem[280] = 144'hfdb4fe6b086001b50cbd0f69f9bb0f3af429;
mem[281] = 144'h0f2cf138079f0e4203b00080f494fa96f68f;
mem[282] = 144'h0bcd013ff2ccf7de0dedf9bef327f7bfff84;
mem[283] = 144'hf0f0f80ff83e033bfaa3fd8d0ddef8950dad;
mem[284] = 144'h04a60eb30586090bf471f7500f7ef41d0d2d;
mem[285] = 144'hfff9fd7af94100960cadfd1cf1000d12fa71;
mem[286] = 144'h00b30a4b0c50050d05b40a53f5e308e9f3f0;
mem[287] = 144'h0ad30b700b8ff6bbf07afc84068cf696ff15;
mem[288] = 144'hf643f70df1500b9ff738f28a0b930cde01ef;
mem[289] = 144'h06cbf9ddfacbfc3b01c90334fda0f6220a20;
mem[290] = 144'h06e500b00a88f20e0814f7d60ee50ec1f696;
mem[291] = 144'hf57af0c2face0da1062ef605f4dff0c90669;
mem[292] = 144'hf2d8f3f204fef54101dc0fe8026d0b55086f;
mem[293] = 144'hf7a40b090a5df78d08d3fdb7fff6fc7106a5;
mem[294] = 144'hf3cef26befa7002ffb8bf9d2f981f3980619;
mem[295] = 144'hfe0e013a002ef79dfcdefe2409aa0b890861;
mem[296] = 144'h0b2cf4930567f3e8069806d20bc70a07f735;
mem[297] = 144'h09790f1d0a05fffdfc360125fb0df91bf3a0;
mem[298] = 144'hfe62f19005e309010ebaf9c203450ad0ff01;
mem[299] = 144'hff9a0406f9ca038bfa33f5d00389efdff95c;
mem[300] = 144'hf70c0d00f932fa4d058af46c014d0657fa50;
mem[301] = 144'h091bf0bffd65051bf38df5480f7309a30077;
mem[302] = 144'h0198ef7ef9dbf5e80a18f16f05d60b92ff2d;
mem[303] = 144'hf1d6f91af532fe1c047304c2fe1900410572;
mem[304] = 144'h04d2f9a7fc4c034cfe8e04650f67fa42f951;
mem[305] = 144'h0e900c8902760bd103aefbdf085008ea0cb8;
mem[306] = 144'h04350f42f0f1073bffac0454f7380b31f6b9;
mem[307] = 144'h079ef23f00590181f650fcff0710f4660110;
mem[308] = 144'h048e0d79fd2d0062f21c01cef7f004aeff4f;
mem[309] = 144'hf26302a9fde207230d220c19f18500d20c22;
mem[310] = 144'h07ddf0f0fdd2fd71f2aff857f4620b1c08c8;
mem[311] = 144'hfbddfbf30492f07c00a0f5a0f638f2adf16c;
mem[312] = 144'h0536009cfb3df8cd06c30ce7fb980ec603e5;
mem[313] = 144'h0f00f012f6a1ffbb00dffe14fae2f42bf416;
mem[314] = 144'hfb71f5a30e940490067c00def48e0343081f;
mem[315] = 144'hfcf4fca40b6f00940dbb01120a35f9840804;
mem[316] = 144'hf770fe9e082c048c0cc0077af28f03ecf489;
mem[317] = 144'h0bd8f478f5bb0c76f747f6f803d0f543f8cc;
mem[318] = 144'hfb5ef61cffc0f93a06db066e0dc6f237f11f;
mem[319] = 144'h0b4e082d00410e0ff27ffa260bf4f73704e4;
mem[320] = 144'hf892f6dcfc210733f9a1ff880ebaf872f256;
mem[321] = 144'h02790761f86a081cf719ff2afbb6f304f5ed;
mem[322] = 144'h025a03f20e8608c90733f9790e1bf0230087;
mem[323] = 144'h001e02cb0f8b0fc6f776f82af872fe290c01;
mem[324] = 144'h08aa03050c150961040e0e30f5de0a2ef526;
mem[325] = 144'hff87f793fe32fe76f1140adc09cd03c8f564;
mem[326] = 144'h0f16fd17f774f6ca066a03de0254f21df46f;
mem[327] = 144'h0a5802930a85056fff6cf24e081c042ffb0b;
mem[328] = 144'h0596efb2f4700121f784fef809b30d4e0de0;
mem[329] = 144'hfb65044906c0f7b90b16f4aaf58ef9490218;
mem[330] = 144'h0998077e05f5fca30aa80413fd91023c025c;
mem[331] = 144'hf1b9f3970c02fa660c44f7f6f590f5b20022;
mem[332] = 144'hf006ef360976f5c404970a72f15defaa040d;
mem[333] = 144'hfaeb0be30468072c0190f93afe1bf8b5fe64;
mem[334] = 144'h008e07e105def29d0867084ff411fd8defe9;
mem[335] = 144'h0287f583f44c05200e99ffe0fb6e097df060;
mem[336] = 144'h09bef58cf1f30ed602a2f2e50f860c1e01b9;
mem[337] = 144'h0637f1eff2a6f49d0e11fa68015dfbcafc2b;
mem[338] = 144'h0903fcd40ebbf857fbef0a910647f54e0db3;
mem[339] = 144'h050802000a4c0dd7f0780855f0fc0c98095a;
mem[340] = 144'h0a79ff39fb1705c00bd1fd6a00ffff39f2e9;
mem[341] = 144'hfd460a500949f69a016bfb4b0ab40b1bf871;
mem[342] = 144'h0c8806330cb801a8fc7dfdf106230f250a00;
mem[343] = 144'h07a0096cf7f1f11ef68af60508cdfb72fc7a;
mem[344] = 144'hfcc206e6fe5cf9def77cfca0fe2307f6fe8f;
mem[345] = 144'h0450ffda02110ec40d3506e7f42000b00f0e;
mem[346] = 144'hfe5c0a7c05f2fbb6098dfd35fb9cf7e5039a;
mem[347] = 144'h065d0be0f0f8f080ffe20d2cfb3cf84a078b;
mem[348] = 144'hf34df2f7059e0d6afe83fbc50de8f17eefdd;
mem[349] = 144'h0d750980f9060b5cf2630f88f79bfb8b0096;
mem[350] = 144'hfb7a097b02710e9104680a2bf15302e2f356;
mem[351] = 144'h062e0b84fc54f114000a0051f3280e89f02f;
mem[352] = 144'h0ea30537f8da0be6fbddf225f529fa34005e;
mem[353] = 144'hf2d7ff35ff5af79d0172f5a90e200b4907a2;
mem[354] = 144'hefcc0788f3b40452f4f30447fcc303bafb7e;
mem[355] = 144'h0c900c99f4e50578f15df398f35b0bb000b5;
mem[356] = 144'h00120d86fc45f8c300250182f0aa04f307c6;
mem[357] = 144'hf7470631f011f616f162f74f042b09f10f1b;
mem[358] = 144'hf484f101fb4d0dd00551f31bf58808cefae4;
mem[359] = 144'h0c300aadfd24fc34f7820c3305dcfc700a60;
mem[360] = 144'h0e80facef486f826fe16f50afc72f8e3f657;
mem[361] = 144'h0a860eac0bf903c1f4b60f790840ff4503c8;
mem[362] = 144'hef860ce304f70246fb000e76f079f9dc09f3;
mem[363] = 144'h0182fc810e080c2ff5dcf86c07900bda073b;
mem[364] = 144'h0c94fd76fae5ff4ef1a6fbe3feaef726f9e1;
mem[365] = 144'h0c43f0cef38bff6007d7fcc8ffb30c830252;
mem[366] = 144'h04460b6507e20095f3590f400e26f432f373;
mem[367] = 144'hf71602e3fc5a0f6708eaf3320e1af913fdca;
mem[368] = 144'h04ecf7cf0e52f755f83fefd80b97003d0512;
mem[369] = 144'hf026fee4f07dfaaeff00085ff0f109760fca;
mem[370] = 144'h0daf00240f9bfc1cfef9f574008500fd0837;
mem[371] = 144'h0cb70f560f76f73bfc91056ef7f3f141f561;
mem[372] = 144'h0dda065f0f9bf1f5fb4f05e2f009fe1d0207;
mem[373] = 144'hf3bb058c04c80b31ff780c2608f4faf403b4;
mem[374] = 144'hf22cf330f81e04480b4af93308eafa7df9f5;
mem[375] = 144'hf9260551fc76f1f60ee40a8a0ab60b32f462;
mem[376] = 144'h040dfa5f06f5f5bc0223f972fad80e970f8b;
mem[377] = 144'h00230626ffb0ff7df917f0b80cc3fb3ff676;
mem[378] = 144'h03a5fa08f636ff0d039b01540c420163f7b8;
mem[379] = 144'hf7fd01410c830f160dccf4fc0871fdc001c9;
mem[380] = 144'h00bcfb7ff99ef35204c0fab10e91fd000a73;
mem[381] = 144'h080905e5025af2d7092c0e66facbf40af142;
mem[382] = 144'hf8380377f5e30c8704bcf3f20dbffa4604d0;
mem[383] = 144'h02b00e100d230ab900a2feac013af0ebfe64;
mem[384] = 144'h0627f02bf3190dbef1e80ac103e60ace0c37;
mem[385] = 144'h0657f1da0f6308f20870f2540f6efdabf71b;
mem[386] = 144'h0c6c058df4140f95f3a50c90efcbfba009b3;
mem[387] = 144'hf094fdcf0ca8fc600d9ef7fd032a0219f733;
mem[388] = 144'h0bc5f5f4f6b00981f9aa08800af2f993faaa;
mem[389] = 144'h0cdd08affa2a06870386f2e309ca02c9f88f;
mem[390] = 144'hfd77ff2df38bfc8005b5f5ebfa860a54f1bd;
mem[391] = 144'hf36809c8f8acf17fefdbf611f07ffcebfdce;
mem[392] = 144'hf438f4abf6a7f255052ff4b401fb0ae4fbe6;
mem[393] = 144'hf8b209dc0f1a0ccc089a04b907e60489f5c6;
mem[394] = 144'hf14f0568090305affdc7014b03b7f3abf6d2;
mem[395] = 144'hfe750038025afe76f75001970eb0fb3cf244;
mem[396] = 144'hfc43f5530a9605b40e7bf3dc007ff2a30a4c;
mem[397] = 144'h08aef9d107000c35faaef7df07ff085f0cff;
mem[398] = 144'hfae50ea70447eff3f923012305ae03adf0b7;
mem[399] = 144'h0f1a0052011efc1ef5730aabfef4fa6bfac9;
mem[400] = 144'hf4f6f1feff480c2c028bf6df056af2fb0772;
mem[401] = 144'h0d8ef39a00fa01ddf8670bea02cf0598f9e4;
mem[402] = 144'h0b650add05140d16f4fafdc3f6b0fe65f5c2;
mem[403] = 144'hf94f02220bb80544f396056f009703b4f7fd;
mem[404] = 144'h018ff8f9fd84ff5809cdf3840bf1f672f14d;
mem[405] = 144'hf49a014bf917036206e8f45205f3fc800a04;
mem[406] = 144'hf603f77607740de8f7a9f5b002bf03ca0923;
mem[407] = 144'h0a41009a0bcbfe4bf932f9d700bef06904e2;
mem[408] = 144'hfeb9029cf67d0198046f0d9af158fad3f6cc;
mem[409] = 144'hf72bf113fbadfcaaf662fb5905f506c70411;
mem[410] = 144'h0590f004f1ae0794f5d606ed06a9018af571;
mem[411] = 144'hfc820dd8f27800270f1cf11f0bc8fec10058;
mem[412] = 144'hfc59ff450c1400cbf4f80b3b0a220f9afb7a;
mem[413] = 144'h01a301480e25f39a0581fca1f43c0e120253;
mem[414] = 144'h0074faeeff81ff2906b3093d07c4f02f06a2;
mem[415] = 144'hf919f31c0816f5f50b5efdf1fcb3f3b1f144;
mem[416] = 144'hf40501a703d7f3ce041ffed001b3040dff0c;
mem[417] = 144'h0584f0200e1bfe3407bdf07e01cc00cff1f4;
mem[418] = 144'hfaa30451fc87030908b904710a3d090af649;
mem[419] = 144'h057a066409f80c50f770fc5c04260a9ff328;
mem[420] = 144'h0733f4700b99fdf70dc10b9007a6fed70672;
mem[421] = 144'hf765fd700908faf30999fc8f0605f727096e;
mem[422] = 144'h05bd07e5fc15f05ff45a03610fb603e109de;
mem[423] = 144'hfe0f0970fe1d0c58f6e0f6b905f3ffac048b;
mem[424] = 144'hff220c54f3f7f4f5f82bf0ddfdcc05c70f5f;
mem[425] = 144'h09f506ac03cdf75d0b8cfdd2053ff45dfac4;
mem[426] = 144'h0fdb0241fb1ef76602c5039e0e4609090391;
mem[427] = 144'hffc10448f94df66f05adfda3f7bcf7610051;
mem[428] = 144'h040eff6909cefe2f02a9f64af454f90ef6eb;
mem[429] = 144'hf06ffe2905ecfbdeff8ef6dc0b440f9c0dfd;
mem[430] = 144'h0f32f631f84ef4850e1b05030632f5c4fcbf;
mem[431] = 144'h02f2fc35f5cafcee0e01fb9103de00a7f690;
mem[432] = 144'h0fcf048f004cfeef0185f382f40b0be5017f;
mem[433] = 144'hf55e01cb0aa304a9f1fdfd9401070efb06da;
mem[434] = 144'h0f64f9cc0cb3f01ff9c705eefab0f5e6fcfd;
mem[435] = 144'h05e10e3cf2a1033bf41407fb0a91029dfd73;
mem[436] = 144'hf5a90234040d0a7c04bbfed5ff2207580325;
mem[437] = 144'hf29a0989f4c9f14ef55cf72ef9dfff340351;
mem[438] = 144'hf074080e041501ce0ac507cfff68f2620d6b;
mem[439] = 144'h035402b3f64af7f200e704c30ebdf5300046;
mem[440] = 144'h0309064df34d0b91ef2ef6cf054d05750513;
mem[441] = 144'h01600e88f5a30988fbb4037dff2009df0a25;
mem[442] = 144'h0bcbf10905a60996fe66f5b2fb6feff5009c;
mem[443] = 144'hf5f8fe82f7da00fdf118fc9c093b03d205da;
mem[444] = 144'hf3ed07800d7ff372fd3df60df2770d02fd8a;
mem[445] = 144'h05f001670d72061508c40899f46cfed30db4;
mem[446] = 144'h0ca3fc2cf7f00374f8a5f09efb06f94d0064;
mem[447] = 144'h002ff81bf8a4fd0a0aa00cecefc60cbdefa4;
mem[448] = 144'hff92fd9e0bb9f7550caeff650e02039af0e4;
mem[449] = 144'hf8cef9eb002002b801a5f8e9f9b7fe820c41;
mem[450] = 144'hf3faf8290abe02c00f11ff7906850d7b08d7;
mem[451] = 144'h0b19fe21f04afaebf654fee7f7cefc600f0b;
mem[452] = 144'hf56df69dfac4044209540530f900fa7cf94a;
mem[453] = 144'h03a5fe220445f8960bdff4170ccbf89a0b12;
mem[454] = 144'h05d7fb22f9900da8f54009a9fecffb03ff5e;
mem[455] = 144'h09830417fbd5fdd90932062806400aa90073;
mem[456] = 144'hfb2fff9cf6f6fbc1fbe304e403cefe40f948;
mem[457] = 144'h06180e390f99f32af033f4d3ff32f00b0f3b;
mem[458] = 144'hfa28f99dfce7094ef3b00e98f674015ef200;
mem[459] = 144'hfc240f81fc09ffe8ffd9fb31f742f7740e24;
mem[460] = 144'h012e073604dc0acaf1b10698fe20fd19085e;
mem[461] = 144'h0d75f22af3150108f60d03d0f8cb0b6a0c5e;
mem[462] = 144'hf0edfa030416f40a0ed8f2ac0ca80981f533;
mem[463] = 144'hfeb0ff27fc7ff4d3039bfd4e09c30eadf6cd;
mem[464] = 144'h0eb80988f9f604f10d9d032e0471041300b5;
mem[465] = 144'h0a72fc000754f2eb0505fdab0b4b08ddfdff;
mem[466] = 144'h0578f33e0c530020002f00a0053af7f70660;
mem[467] = 144'h01f506b1fcc90a3cf1ce00f608b300290beb;
mem[468] = 144'h08eefa7bfef4fc710a5607ea0606faeffa62;
mem[469] = 144'h0b8f0d6ff936fed50888fe400293097cf93c;
mem[470] = 144'hfc020f2cf4e0fa2c0354fc190fb9067cf072;
mem[471] = 144'hf850f46b04def35b05a70c400afff423fbe5;
mem[472] = 144'h02490953efe2f8d2f863f7c006d4f9a6fa4f;
mem[473] = 144'hffcc0decfb86f8d30877f3440948fa070380;
mem[474] = 144'hfa9df4d3f44c029e096a07bbf0470c440cb8;
mem[475] = 144'hfe7f0d920b29009b06bb02f20a01080cf26d;
mem[476] = 144'hf7c3fb0f0f31f82b09e9f43005130c4c06f7;
mem[477] = 144'hf25c0f88f2e80caef8dd04c4f6b6efe6f27d;
mem[478] = 144'h0af1f5b90dfaff290e5c05bd0d28fa110c88;
mem[479] = 144'hf8a201ba09470f620599ff28fc9a0985f9bc;
mem[480] = 144'hf9ce0fe4f8ab030802860668f824f154f34e;
mem[481] = 144'h0181f1b5fc08f358f25b0af7f18e0d3c0eed;
mem[482] = 144'hfe7504bbff58fa41f6fd0a1a0f670ba0f8a7;
mem[483] = 144'h084f0a700be5081ff6b70b6af1f00e62f7b1;
mem[484] = 144'hf0020e730f58fc490f7af6620154f26df5bd;
mem[485] = 144'h07a20bb90d0dfb7afbcdfb5f03bcf12ff9b4;
mem[486] = 144'hfb62f2f007c5fa52fb510b6b0506f8920bd1;
mem[487] = 144'h09a1f81af0270e88f9c7f0b3fbccf287fb65;
mem[488] = 144'h0209f8b5070ff260f2daffd508b2f889fb36;
mem[489] = 144'hf12c0250f926f793fe870c3c015602a50596;
mem[490] = 144'h0ab7fff4fb0d0366f7b4023401f30377f219;
mem[491] = 144'hfd4dfa56f910f0f2f7370ae70675fbd0f591;
mem[492] = 144'hfc05fc11084b0536f74a0accfb540e79ff66;
mem[493] = 144'hf31a02b604db0e5a0c9b0dfd0d88059af7e6;
mem[494] = 144'hf1fb0042ffcf07fbfc070655fcb5f674f792;
mem[495] = 144'hf33df61c063605b00092f29c0edff1930602;
mem[496] = 144'h04c8f8def83f0af6f9730b39fb99fdabf9d8;
mem[497] = 144'h058ff986f5dc011903a30f46f28603d2fcfb;
mem[498] = 144'hf8c304b1f741f4ab0afdf710f34afa8f0ef8;
mem[499] = 144'h0c5d0901f9c207b1f9fe0f65f1a50b09fb1b;
mem[500] = 144'hffd60225fa120074ff580af406fef23d0695;
mem[501] = 144'hf18803a50ecff8a2fe0807bd00b6facef4b3;
mem[502] = 144'hf83af87c0529f2240d16f5ae02dffb570de7;
mem[503] = 144'h087cf3a30a730d6afdfaf289f3eef23ffacf;
mem[504] = 144'hf157016cfa54f8bd038dfdad02ceffb8091a;
mem[505] = 144'h0e9400e50e7ffd450ceaf7eb0bd00d6f0269;
mem[506] = 144'hfc36f9cefd7a029af01cf63d095b0c6ffacc;
mem[507] = 144'h0487094bff13fd1e0b79f0f00328fd2ef7e4;
mem[508] = 144'h0a53fdc1089ff1400b0705aaee83f9ec00ab;
mem[509] = 144'hf5edf4a6f4e40669fe64f26a0c820007f5b2;
mem[510] = 144'h05d909fbfea8ffb709930186f3f0f1f00dd2;
mem[511] = 144'h0dc1071a040bf7dbf235f6d5f1130b3f0b9c;
mem[512] = 144'h09fd050cfbc8f002f18cf0d60a01f3b2f8c5;
mem[513] = 144'hfa29f48ff6f4f11408eaff2b0bc20d760e9d;
mem[514] = 144'h0dd80df202450b450ebcf7d5f282f9f6fdc8;
mem[515] = 144'h0941f08c0848f4e5f0d8faf10dc7fa08fed3;
mem[516] = 144'h090c0166f720fb50f04af819f268f6f80ca3;
mem[517] = 144'hf8e7f90cfc7cfc7a0a0e0200f40f034a0528;
mem[518] = 144'hf492febc018a0e1cf795f4ac0b1efa02fe94;
mem[519] = 144'hf385f9d40222065dfa8e020a0b41ffc50183;
mem[520] = 144'h009104d2f50cf21701790e900993f5cff64f;
mem[521] = 144'h0e08ffcef6bcfc73feab02a1f330fbd1f593;
mem[522] = 144'h0ab50e570df2f2ec05e2f911f6de00da0549;
mem[523] = 144'h06e4ef93063f02170a21f77f0430fdd60a46;
mem[524] = 144'hf6880c1b04a6f7caefea07130c7fefcdf4f8;
mem[525] = 144'hff1608fff50bf7ad0c84f3ce09ef08dd0abb;
mem[526] = 144'h0518083b058c023e068bfb830ef30a52efe6;
mem[527] = 144'hfe5206d4f67ff570f70df90b044dfe80fafc;
mem[528] = 144'h098004c3fe690c2cfa25f9a9fdfff4240e76;
mem[529] = 144'h03dc0675086e02640cb5fbfdfa51013e05f0;
mem[530] = 144'h010bf77cf6920dbffd2f00820fddf8380648;
mem[531] = 144'hfaf2f1b102260a2afc39f9a30e40f416fdc0;
mem[532] = 144'h08c1f562ff360c2808b7f6c2fc31f598fed2;
mem[533] = 144'hf683082ffcbcf3640dc7fc8cfe200538f720;
mem[534] = 144'hf96a0c910ae409e60e9d0788f227f839f189;
mem[535] = 144'h0023fd1e0656f1dcf96c0f27f0f40b100062;
mem[536] = 144'hfac3f6d009cc0a4ff8e8f4cc086d01adef8a;
mem[537] = 144'hf95a0b9dfa5cf1cafa1b02e9f63df6a5f9cc;
mem[538] = 144'h0d1b0331f6fd0d09efd0f83df1a4f15afea1;
mem[539] = 144'hfbb1fcd8f1f70af7f34904640208f774ffdf;
mem[540] = 144'h077ff396f28c07ac01cf08c002a7f045003e;
mem[541] = 144'hf39df86e061e083703a80efe01c6f7b8f32b;
mem[542] = 144'hf0280b78f764ff09f41208bffd0006820e2c;
mem[543] = 144'hf2190f82f9f00b31f921fb9ef9b10ccff2ba;
mem[544] = 144'hfd0ff5f4f844f7b70e39fad4f04d0394029a;
mem[545] = 144'hf8c2f4c80756f1e1f926fedefb8af9710b4e;
mem[546] = 144'hf454fe1408ba0051f9ccfc970e8708c60b96;
mem[547] = 144'h0cbd0cd9fe90ff370f2ff159f5750e3efc28;
mem[548] = 144'h006a0257fb99f86df3610e47046bf326f1cf;
mem[549] = 144'hf57d0be408af078ff5c409bc0c090c0fff3c;
mem[550] = 144'h024c07f706a6093f07510251fec009a9f6ef;
mem[551] = 144'hf0bff8a6faa008660dfc0127f62104f4f24d;
mem[552] = 144'hf731095604570891fa3ff5ddf5ad0c3bfbdb;
mem[553] = 144'h00490fb6f41ff87503750628fc8cf0a0fb89;
mem[554] = 144'hfb5a00e1fe0ffb980a04fedb07baf3720ac8;
mem[555] = 144'h0513fdf9f3bafb01fb29f699f16b04ed0493;
mem[556] = 144'hfee2f53df8edf7170d4b0f3c0f3f0c35f629;
mem[557] = 144'h00220680fd040c0c001ef0a1ff2ef610006a;
mem[558] = 144'h08710950f79df634fda7f478f647f5c0f173;
mem[559] = 144'hfada03d2f17406a0fb1ef068f8040a4dfe4a;
mem[560] = 144'hfebef34c04faff75f94402c30ce7f5d4f9d7;
mem[561] = 144'hf1a70222ff43f281f366fa3a0bec0629fc6e;
mem[562] = 144'h0fd7f4870c2bf27b09a5f9dcf8f00c1307ab;
mem[563] = 144'h0f690166f21a04a40e4df26b0a31fa4d0a6e;
mem[564] = 144'hf2d0f7360250f7c5f8c201110d95f493fa28;
mem[565] = 144'h047bf69d04be091ef7bcf041f8f1fda20be7;
mem[566] = 144'h0e65faf8018106a602310f340238052ff54c;
mem[567] = 144'h0e60f35c0e21f1b703010c4f043608e7033f;
mem[568] = 144'hf0dafca3fbfbf3b0f03d00b9f9e3ffa60962;
mem[569] = 144'hf2a80578fd9801d5078201ce0928009af9bc;
mem[570] = 144'h036a037ef50ef650fe140e1cf857fd090ebe;
mem[571] = 144'h014dfe580c48f63a0a6df287fb790191f08e;
mem[572] = 144'hf5260d2807cbf20bfce4041ffc66f874053e;
mem[573] = 144'hfffb0391fa0e011d0e0afe2bfb5a0a96f797;
mem[574] = 144'h0e040ac300fef439097f0d2dfb3cf825f495;
mem[575] = 144'hff060132fcfffb7d06c9f471f504f1d4f1a8;
mem[576] = 144'h0d89fd6b025bfa9ff829f57e001f0159fcff;
mem[577] = 144'h0126027bf0f002fefb94080cfb23f4840fc3;
mem[578] = 144'hfdfdf2360e8df9480702fc160579fd7b0a35;
mem[579] = 144'hfb440e1808cdf85ff6440006f4edfc73084c;
mem[580] = 144'h07680e7a0908f8e400040b7d0bc2fcddfbdc;
mem[581] = 144'hf56005c5fb43015d00360e180c0104e8f867;
mem[582] = 144'h048ff068efce01840b0ef2d1f14af2970cee;
mem[583] = 144'h0e8ef65dfa76fda6f67c082907b90918fbda;
mem[584] = 144'hff0cfd2bef7df139f7a7f1770224018ff05d;
mem[585] = 144'h0afdfae1f287f751fbb60cc1faf008a407e4;
mem[586] = 144'h0bbb05c9fdb70cd509d4017d04b8f5380a94;
mem[587] = 144'h0c9b0a44fe07f7d80298094cf5e30913f36e;
mem[588] = 144'h020b00bff9fc0640f3dcf7bbf4fcef79fd95;
mem[589] = 144'h0ba900c10e740f140be4fcb305fcf930031c;
mem[590] = 144'hfff50d6bf35901b305c0f27bfed901a7f324;
mem[591] = 144'h025c032e0696f00003ecf3fc05c0f8f3004a;
mem[592] = 144'h00ac0cbcfe9f036307f20c1d07a7f8b60103;
mem[593] = 144'h04c403c70fa6f08dfad80ddefc38feb6fa8e;
mem[594] = 144'hf3faf75a01cff59ff1220f940dcffba0f795;
mem[595] = 144'hf44a0719f65ef9f8fa350225033a0d3df244;
mem[596] = 144'hfc4a0b5302ce0b090bce0c35f0290c1804c5;
mem[597] = 144'h0314f6d901dc05cef7160d04fb43fecefc17;
mem[598] = 144'hfd5efd0a0cf104c7075f034eef74017b0194;
mem[599] = 144'h0357f30305d208baf1dcf87b011df683062c;
mem[600] = 144'hffe30378f62d060c0ccc089809d6f9940391;
mem[601] = 144'h0f76066af22e0685fdef0e8af6620cc4f53c;
mem[602] = 144'hf196028800b207ac06df0284efb00e1bfda1;
mem[603] = 144'hf22dfa3afe4df3760cb804c30bc4fd3e0242;
mem[604] = 144'hfccd0075f9a40149f315f546fa22fce80cc9;
mem[605] = 144'hf56a001309cb0343f057f914fff4f65ff172;
mem[606] = 144'hff2b04b00ca40a600c5e0f9c0ce4f9310a52;
mem[607] = 144'hfbb30851f40e0268fa0808070fb9fba80d10;
mem[608] = 144'hff120d32f728f0510d8c0f6a078e07ea0e44;
mem[609] = 144'h06640e4503e603b1049cf191022201c0f7b5;
mem[610] = 144'hf0090cdaf5380cc20ad2fa5ef2eaf16efcc2;
mem[611] = 144'hf75e0b38f93cfae501d7fea6f9f9f835fb62;
mem[612] = 144'hf5b804980b4902280da2f0bdff2705a6fee1;
mem[613] = 144'h00e2f13c05ff057efd30f9d208580a27f3f7;
mem[614] = 144'hf755f324fdc700fd0f2af0fff31ff8590a4f;
mem[615] = 144'h01620dc8f8dc0738025bfa4e08baf9ecfd68;
mem[616] = 144'hfacb099bf8b106c10ed706ed0aaf07e30bc0;
mem[617] = 144'h08d20ce800410a0b0b0f057ff1fff664f052;
mem[618] = 144'hfa68fde4f0a50bbdf47e0f120aee096303d6;
mem[619] = 144'h03710ab4020d0a8806ae0b96f2890947f61b;
mem[620] = 144'hf18df870f49ef29d01860e5b048bfa0503cb;
mem[621] = 144'hf792f3a8f9fcf8eaf59df51ef404f4d2f05e;
mem[622] = 144'hf33e090805510d10f3dcfdfa0f29f1bf0acd;
mem[623] = 144'hfbabfc760a49fbdff72605e709290691fd3c;
mem[624] = 144'hf6300008fdf3f2e8f47bf22bf35af2eefd7c;
mem[625] = 144'h070100ed080202dc0a32f3de0d5f02a60406;
mem[626] = 144'h03f4f2affd26fc6efc94f1c30b550db5effe;
mem[627] = 144'hf6cc0699f78c081a04bf0fe4f7780f7a0120;
mem[628] = 144'h078b0d1df13b08bbf5ba07fcf9bd048f0214;
mem[629] = 144'hff2c0b6ff1daf11c05dd0544fbc7f10407fb;
mem[630] = 144'hf1fb09ae06e00072fbb4011af6ff0dd70326;
mem[631] = 144'hf1cbfebf04e3fb3304c4ff64f9880dbe0c60;
mem[632] = 144'h074afe680412f254f6010a950810068dfc28;
mem[633] = 144'h0275f1f40c83fdf201070833f51f09f2fa87;
mem[634] = 144'h0474fca70573fdf206b9f9caf3b308fa01b6;
mem[635] = 144'hfc4ff924f80c088105720686056cfdb8f1d9;
mem[636] = 144'h0cc1fc9804c3f6680a09fe81f2a3fc51f915;
mem[637] = 144'h08fe07dffe7bfd58fbe4fc57f80d07970263;
mem[638] = 144'hfb680aeef1cef60af02f0adafda90a95f625;
mem[639] = 144'h05400f4d0136f74301460236fdcef93c07bb;
mem[640] = 144'hfec4f5caf54bfdc308040e1d0ef8016f0819;
mem[641] = 144'h032ef48ff0020ba50185007a0d87f990fd61;
mem[642] = 144'hf0e5fd7801cefd24071c055f0d30fb2f07f5;
mem[643] = 144'hfdd0f456f228f08cf50b021d0767f3420a93;
mem[644] = 144'hf67ef4c80e36f32808f5f5fe02cdf2edf5e7;
mem[645] = 144'h0a9d00b6f7df06c9f29ff06df5050aabf94a;
mem[646] = 144'h0f760e95f29df9dd0c69091c0603f8f0044f;
mem[647] = 144'h0c79ff2afcfbf1ac0c67feae0422fc15f03b;
mem[648] = 144'h0a180d30f82307bbf716f494f376fbe6f09a;
mem[649] = 144'h0a10001ef40309920ad9fd600a4ff482fc0e;
mem[650] = 144'h06290158fb350926ff680caef832f715f7f1;
mem[651] = 144'hfbf2f82809acf0460b6f0c0ff80b01fc0218;
mem[652] = 144'h0f6504960c6fffeaf22e01d2f3820e6f03aa;
mem[653] = 144'hf03df6160df7f4e90597f4d500ebf1d7fdcd;
mem[654] = 144'h085a07c707ff010df669fb5bfa0cf712f16e;
mem[655] = 144'hf5b90bf0f011fbcff7aa082bf6df0df4fff4;
mem[656] = 144'hf82bfed30decfeafff1efeabfebdf3340544;
mem[657] = 144'hfba8fb95fccdf587079f00c20210f2f0fd65;
mem[658] = 144'hf74e0098efe5ef480044f9e8f4ac06f4000e;
mem[659] = 144'h07160e990de5fcecf74302d508eb045df051;
mem[660] = 144'h056dfc9dfe7904aaf73d0b75fbd50a460a95;
mem[661] = 144'h0cc00146f67c0d8ef8190b6afc77f92d0f4d;
mem[662] = 144'hf66209d00b98fcc4082204cd0dedfc5402fe;
mem[663] = 144'hfba20dd00920f38e06ef0e81fe8c02af0dc6;
mem[664] = 144'hf1150ef60d48f72503a5ff5207f5f9cf091d;
mem[665] = 144'h08e9f685017a03260a3701ebffa5f77e0e9e;
mem[666] = 144'h0be9f65808faf3f9069afc4a05590caaf8b9;
mem[667] = 144'h0955fb56043af4e3f8c200e3fa0dfc3afd43;
mem[668] = 144'hf89ef903f732fc4c046709aef994f696f005;
mem[669] = 144'hf5cf081c0b6b034af42d091cef480cbf0293;
mem[670] = 144'h09c1f3940167fd95f5f30f2ff89ffbbafbae;
mem[671] = 144'h0beaf8c50b6c02a104230cf50f1101d0f9d0;
mem[672] = 144'hfa9bf93bff89fa38fdabf3e00cef0c03f054;
mem[673] = 144'hf0cc068ff040fbe8f5c708880bd4f86007cf;
mem[674] = 144'h06360a36f36b029802bff11301860026f0d4;
mem[675] = 144'h0e5efe7df88b00360be3f7d7f36bfb0afbf4;
mem[676] = 144'h09f4098b0774f98a00c50d1afc800a1b027b;
mem[677] = 144'h0af1fc37f8d30ca601a50146f0f90552fb60;
mem[678] = 144'h00c806f00473f920021afa360d0c08650b56;
mem[679] = 144'h0471042fefdc0d4c02500e2e0a7cf6c80122;
mem[680] = 144'h01200909fb4e09870c24fc5807fef13ef9c0;
mem[681] = 144'hf4ca056cf28fff21f90df1280c9b0314f3fd;
mem[682] = 144'hf8d2fdf3fad50ed3fc0b03b50998096c0dc6;
mem[683] = 144'hf684f635f6aef55efab9f12c07db0956f800;
mem[684] = 144'h0fdc0f7cefddf02afb51089ef7ee090b0c11;
mem[685] = 144'hf3ccff800a88f311003c08c3fcee0254f199;
mem[686] = 144'hfb9105c10f2ffde5fc4c0da1f24606b808c5;
mem[687] = 144'hfa4bf265040806840d540705f70afdc807d3;
mem[688] = 144'hf4d9fc940398f6d303e2ff37f2a902e1f833;
mem[689] = 144'h049cf1d9fca3f0f9f7dff203f59ff13b09e2;
mem[690] = 144'h0c1309e2f02307c00371f0c20c42fd20f637;
mem[691] = 144'hff5004a4057103920fad098f00daf7240b50;
mem[692] = 144'hf7e6fa1bfd6d0452fcd70d7bf4100352f0a6;
mem[693] = 144'hf57902f0f7e0f8c70ef5fbfdf7c504f50e33;
mem[694] = 144'hf20cf146ffb5fa08f379f302031afe97f232;
mem[695] = 144'h0d6909980860f79cf80e0392f044f83f059e;
mem[696] = 144'hf0f303b6f103f481fb540eea0c3fff9df8cb;
mem[697] = 144'hfa9af7fa0ba30b4800e1f2b6f78b06ecfadf;
mem[698] = 144'hfaee06b901b9f9c7fce1094df86908490ca4;
mem[699] = 144'h0eecffecf599f0c8008df38e0f6a0ac6f790;
mem[700] = 144'h01720742fe25f34af878f91c01c1f4dbfa60;
mem[701] = 144'h0b58fd7502920857fdc8fd66f1f1fbc80787;
mem[702] = 144'hf19d0a66f71707be06670ac6fb7c013e026d;
mem[703] = 144'hff5b08b201a009f404f300d9fd9df71b0809;
mem[704] = 144'h07bbf60b05bd055ef49401f30517fe98fba1;
mem[705] = 144'hf0b9095bf72ef982057bfc47032df4cef81d;
mem[706] = 144'h067ffdd4f6250e1ff1f0fe8a0b000e9e05f9;
mem[707] = 144'hf0e80e7df107fbcbf8baff4d0c49f1f2f0d5;
mem[708] = 144'hf49ff6e8fb7bf0c1001ffef2fd3ef1d2ffa8;
mem[709] = 144'h0df403f9f05405440fc6025cf6d703a6f623;
mem[710] = 144'h0a47fa1602cef82b0b2bf312ff2b03e2068b;
mem[711] = 144'h0242fbc9f5b1080d06440d89f87e053009e4;
mem[712] = 144'hffae052d011cf055fe7ff44cfe65f6bb0258;
mem[713] = 144'hfc700e49f6650654095d09420868f84e0f49;
mem[714] = 144'hf90ff58df58af511047cf86008630859f984;
mem[715] = 144'hf2560e33f4640771fe1bf9340f72090ff675;
mem[716] = 144'h0b2bf88ffd25f4dbf3b70b1c0311f8b3fa17;
mem[717] = 144'h020b00a70e82f62d09c60b99008b0c0ffe31;
mem[718] = 144'hfdce0f0306da0db309980581f4f5092a0c07;
mem[719] = 144'hf030f08c079b05940043f476f2d2eff9f526;
mem[720] = 144'hfae00297f04afba1f911fbaff6ce07f2f3ed;
mem[721] = 144'hfb0809c9fbf5f02ef0c80bdaffd3faa9078f;
mem[722] = 144'h0b3b0b5ef4c00759fb0ef53f0041f949f06e;
mem[723] = 144'hf81ff7460e43f3bef196f463f668f770f4b5;
mem[724] = 144'h0751f59ffc30ff730cc4fc460e660d7a0901;
mem[725] = 144'h0970f5c4fd4e0867f76efa6b02c20967fbd9;
mem[726] = 144'h0a3300f9f786047f0095fba1fbe20a3c0cde;
mem[727] = 144'hf41ffcaef1b7f3910401014af5b60d21f0f0;
mem[728] = 144'h0a9a0d420f1dfcb7f711f777fa9e08630399;
mem[729] = 144'hfb000642f0bef8dcff0809af0f6af71f0f4d;
mem[730] = 144'h024e0466037ff458ffd2fa9cf53bf16303da;
mem[731] = 144'h0db9f8fb07a5f6660a33fa730584094ef33e;
mem[732] = 144'h01b5f99df8b3f075f5350afff66206c0f225;
mem[733] = 144'h0d9dff140f85fe3bf0e40a8905f8f9cefd11;
mem[734] = 144'hf652f0adfde30fd0011e09a00846fd74f8db;
mem[735] = 144'h0a580b64083f0fc8f62f091ff082047603e0;
mem[736] = 144'h0a8c0650f2cff9510b01f6a90c7d0d490cff;
mem[737] = 144'h0ba7f51d037f095c0c8e0f890026fad0f1dc;
mem[738] = 144'h06b4089a0675f53e0ee8f0d60d28041f078e;
mem[739] = 144'hf48805d4f1d6faf80c35fde900c20ab80c36;
mem[740] = 144'h080d0817074c0ed7f44c0ae9fccef7c3f1bf;
mem[741] = 144'hfe780df5fba20faa0ba4f35d0169089df6e0;
mem[742] = 144'h0f86fd6ef1ddf5b505f108b9fb16f8a80d7a;
mem[743] = 144'hf61af61807b40cd6053207da0f0f021ef355;
mem[744] = 144'h064a0efc00a2f3030b9b07470359f28af328;
mem[745] = 144'h03330cdaf72307c50513062f0036f1cef545;
mem[746] = 144'h09870a38f062fe28fb0bf782fe07063afe91;
mem[747] = 144'h069e0d13065f0a4ff645f864057f03cd0ce9;
mem[748] = 144'h003704e5fe6ff109fd2302a2fef4fb0c0cd2;
mem[749] = 144'hfaf406dff6a7ff01f5da069afe4703870cb8;
mem[750] = 144'hf266f5e8f2b9fdf9038c095409faf419001d;
mem[751] = 144'h051a0903f047fe51f3410ea9faddf4eb0c5a;
mem[752] = 144'hfa94fd700acd0b470a150b230ee3f306fb23;
mem[753] = 144'hf1a8f6bf0c18fded0abcfe64fbb0f7110c48;
mem[754] = 144'h0bad094e06a608da061808b7f8750c2600eb;
mem[755] = 144'h06410978f580029f029ff02b0348f2caff5e;
mem[756] = 144'hfd2cf94504c80494f018f372f451fea7ff1b;
mem[757] = 144'hf28b0ed90415f3e20560039209fd05daf09e;
mem[758] = 144'h019701b2fe570a6d0b1f004ef82b0241fb27;
mem[759] = 144'hf2e0fe74053f00dbf6ec0938fc790efcefdd;
mem[760] = 144'h0fbd05a8f38cf4fa0c5cf905fc28f8fe0387;
mem[761] = 144'h08ed09aef72a01e3fa320efbf357f01f08f8;
mem[762] = 144'hf12a0001f45d02e3f575f9b10d3509cf0b63;
mem[763] = 144'hfd4300a809ccf96a0b65f655fba1fea6029c;
mem[764] = 144'h039bfc39f08e0a8404080cfc0f630b2209d2;
mem[765] = 144'hfaa1f77c026f048e09810d28ffeff5ea0136;
mem[766] = 144'h0966f49306bafdd3f2ac0d79f0b308dafac5;
mem[767] = 144'hfb71f0db0236f88604aa061707740e800e42;
mem[768] = 144'hfe530258034cff64fe99fd49f4ca0775066b;
mem[769] = 144'h03b60ac5f085fc73060509fcf59807a90e03;
mem[770] = 144'h0edaf51907dd0cc3fa4bf42704ea08230bb6;
mem[771] = 144'h0056fed004b40664fe2305170a80faf803a2;
mem[772] = 144'h0c1b0923f15ef9bfff23ff2f0ea501d40dc6;
mem[773] = 144'hf95907350162fe2a0021f01404ac0ea8f655;
mem[774] = 144'hff920e400c560da2f75002170287057d04a3;
mem[775] = 144'hf27c083709acfcaf0b420b93f071fcad0205;
mem[776] = 144'h02d60f3cf30300190981f45bfd130107f91c;
mem[777] = 144'hfc3a0911fd3306b707ad0c97f3a8f641f746;
mem[778] = 144'hfdb0fb20f452f9d4fcb8f163f54aff27feca;
mem[779] = 144'h0ca0f09b0f53f9c3fae5fdaf067fefebf316;
mem[780] = 144'hf524fd70082f0d690d87f1b30f400d12f487;
mem[781] = 144'hfdb7f157ef0bfa61f981f836f02dfdf10d4c;
mem[782] = 144'hf76401d209a1fff1faf3f8b60d210e9005d6;
mem[783] = 144'hf4ca0976f028f019f8d2f0b60a52fdebfa5e;
mem[784] = 144'hfe4ef72d0ea60b29fbacff37f22d03a9f6e9;
mem[785] = 144'hfca0fc35068afdbff0d7f232f00a0a08fd14;
mem[786] = 144'h0e7705f10e4b03230f9800a80ee7f43cf9e9;
mem[787] = 144'h0a38f1b8fc45f9a2fc1d0eea024403dc08ff;
mem[788] = 144'hfd680c55fa04f3580c14f4e7f5cc0f3afa6c;
mem[789] = 144'hff5406be08c50dcc00c90ce00bcff099f96f;
mem[790] = 144'h02bb08b3fce80bc0fa950c14f53bffd50674;
mem[791] = 144'h0828001ffe9ef73ffb3d00ab0580f7bffc94;
mem[792] = 144'hf65bf1d1f7bcf5570c27f553fc95f4f90883;
mem[793] = 144'hf9b0f372f60009e809e70105f5a1f64201e3;
mem[794] = 144'hfca0f790f518feb401c3f0a8fcba07b8f741;
mem[795] = 144'hfe6bfe87f7670beef7db03e400770708f90e;
mem[796] = 144'h0d46fa5efdcff59bfbe4ff3b01e0f6550f2a;
mem[797] = 144'h077d0781fbe1faf8f5b1f36c00f7f9ad0e43;
mem[798] = 144'hf12d0ed8fc85f9c2fe75f314f2dd0da1f8fb;
mem[799] = 144'h0e5b0d0606910a5b03edfdd6fa06f533f8ea;
mem[800] = 144'hfb0cf24a0ab703f40a5cf39ff7d0f823fa4d;
mem[801] = 144'h0bbaf38dfed80809fe820886f2fdf6570be0;
mem[802] = 144'hfa85013bfe490e1dfede01f20e89fab10c78;
mem[803] = 144'hfb4df4570fc308ef0d2f06f0fb4505ed004e;
mem[804] = 144'h0c6c054b0702f750f579fa9b0ae3f8c10c89;
mem[805] = 144'h0bea01d4fbfaf228021a01f5f1b6f9cd08cf;
mem[806] = 144'hf4f6f94306e609540343f2d605b30d37f783;
mem[807] = 144'hf3b4fe69ffe40e72f6c1f689fe3af41f0d34;
mem[808] = 144'hf03a0923fca60f16efdfff27fbfff02ef737;
mem[809] = 144'h0a030a05f368fc250d7cfb4f073d04a0f072;
mem[810] = 144'hf6f7f10b01df0a2bf19808e2040ffa9cff0a;
mem[811] = 144'h0975f8b80123ff76078cfbc7fa240981fa71;
mem[812] = 144'h0bb7034500710c23ffe2f5440ae404d5f56c;
mem[813] = 144'h0632fdf0f955f6540b890c4ef2af0aecf609;
mem[814] = 144'hfeab0a8f0d2002430936041cfa910d88f350;
mem[815] = 144'hf6d00d00f9fb020ef48207ea007dfd75f6f8;
mem[816] = 144'hf050fd0607d000f7f093fad6fd88f14507b6;
mem[817] = 144'hf68a0c470b56f862f56b061bfbebf167f21c;
mem[818] = 144'hf3500308f7a80551fdec007d004b01a7f69f;
mem[819] = 144'hf0f1fc17f817f2f8f888fb8deff70de206ab;
mem[820] = 144'hf61bf1ba087bf058f401035dfc5f09d7fa59;
mem[821] = 144'h0e5bf5a30ccffa45030604d00953ffc1fad9;
mem[822] = 144'hf66e0b21f48bf170f93dfb70f3070c360868;
mem[823] = 144'h0afa0899f5de04d4ff6602700ca9f31a0658;
mem[824] = 144'h003c031b080e0e14f12ef73df1470930ffc1;
mem[825] = 144'hfaa4f3d601cb08ce03c90c50fc440af8036a;
mem[826] = 144'hf6d00a93efc7f8cc04000b38ef2fff6a00e3;
mem[827] = 144'hfca3f3b2f08dfa6afb38fd1e0af00a240db3;
mem[828] = 144'h0bde0455020ef40f0858fd4bfec20addfba5;
mem[829] = 144'h098a0445054ef06ef2e9f0b4026efd310074;
mem[830] = 144'h036af75ff90506500ad80936fbb1fa0c0a89;
mem[831] = 144'h0b480c53f808f4a8f8f005b7ff52090efaf1;
mem[832] = 144'hf7e1fecef06d09a303780895f23b04c3f14e;
mem[833] = 144'h0aa90ee5f551024c0473f3fcfd1e067508fb;
mem[834] = 144'h0217fbff03ed0761f7e5f62af45b024cf491;
mem[835] = 144'hfe920bb705c1f5500f320550f9330cd6f778;
mem[836] = 144'hfccf0b240043f9b80949f5700f81f411ff93;
mem[837] = 144'h0f42fc3d0aa0f6590f11fd36f53e0501094e;
mem[838] = 144'hf58b0f74f83ff651fb6309d6f6c60f38ff86;
mem[839] = 144'hf150f69807a2f2320769fa70fd44f4e7f413;
mem[840] = 144'h0c3ef5a8fb90ff57012ff3bd0742f4d8068a;
mem[841] = 144'hf95902abef9d0646f445f2baf0950103fda0;
mem[842] = 144'hffd1fae5073a089af88505b801080882f2fa;
mem[843] = 144'h0212f08cf165fd1efb60ffc3f1b70976f443;
mem[844] = 144'h0a58f38107a209fdfbecf3d3f8030f7dfe4c;
mem[845] = 144'hfaf1fbbb0dcefdfef70f0ee6f3170923fb5f;
mem[846] = 144'hf715f0f30b94f8d104170498f8730f49fdde;
mem[847] = 144'h019c0262f1d700370bff0b800c390a5df5e0;
mem[848] = 144'hfdc60b8b02ff0e8f03f002cc0d8afb4b059f;
mem[849] = 144'h010001e3f516fc95f55d01210190045705b0;
mem[850] = 144'h05820534086c0238f98ef5d600bdfd37f8d4;
mem[851] = 144'h0472fbb4098bf506002af45c0c3bfa1cfcec;
mem[852] = 144'h0ab60899fa0df0a4f6890982ff26007ff6a3;
mem[853] = 144'h0dcf0169ff42fd8bfa2cf2910cdcf2820dff;
mem[854] = 144'h0ecf080dfd16f88b0e9c0276fea4fdba0eff;
mem[855] = 144'hfa8bfb07eff502f10383fea3f6ec040602ae;
mem[856] = 144'h043200b90393f750fee9fc6b076a02bffab3;
mem[857] = 144'hf71d0d7bf5b40e3d0a23fcfcf60bfd1f0d70;
mem[858] = 144'h0cc00263f815fec1fb0bfaa10c8d0ba9f9f7;
mem[859] = 144'h0a2cf7e90c4ff908f82d0b2ef858fcde0cae;
mem[860] = 144'hf24f020bfd2afaac09aaf8710944015ffc3b;
mem[861] = 144'hfb91fa0d08ae04690d5f0d7107eaf715f514;
mem[862] = 144'hf0f6f3cc0271f515fab901bcf481f712f94a;
mem[863] = 144'hf6cf02a9f2b203f0022dfc8bf8caf3180e69;
mem[864] = 144'h09e7f7560bc1f092f8b90df7fb11fa3dfb05;
mem[865] = 144'hf4f4f97b0d56f5550005fda30bcb01390a37;
mem[866] = 144'h0796fd480f44fc19ffc308c5f3f8f41ffb5a;
mem[867] = 144'hf75bfe8cf33905b30e30f22e00f508600774;
mem[868] = 144'hf3b60f2f0b75012af8d5f30af235fee6f16b;
mem[869] = 144'hfd5e0635f590f87af64ef13e03c2ffd4f19b;
mem[870] = 144'hf04a0220fdaaf686fa6bffd2f1fa048cf55c;
mem[871] = 144'hff3f014e09c1fd0dfe50f02d006d09efffd1;
mem[872] = 144'hf775f054ffc8095cf06efca306bdffd70cbe;
mem[873] = 144'hfa950fc9050ffa57fc1a06dafa55f7440ec6;
mem[874] = 144'h04d20d12f55efd340e010550fd08082904f7;
mem[875] = 144'h01760afffdfbfc9c0293f909f779f8b70de9;
mem[876] = 144'h0dc8080a08c503d30592fad90536fc0ff6d2;
mem[877] = 144'h040bfaf8f9f808d10b330634f295f704fb88;
mem[878] = 144'h0acd0fcd058bfb53f0560f87f47cf7a5f8c0;
mem[879] = 144'hfb750ced06ae0c0f0bd105d9097c05e707a0;
mem[880] = 144'h0e18fe8cfd6df52df3a9f266f724fe7b090c;
mem[881] = 144'hf70cfdd40c9af52d0dbcf568fbbe05ec0313;
mem[882] = 144'h0aacf232f36d000a0ec70dc9f0befa4cfb13;
mem[883] = 144'hf707f047f2d0fdd80e8a0fc70bbe02f80539;
mem[884] = 144'h04bb0274f27a0dac08fdfb0e03a6f5c50de6;
mem[885] = 144'h0ba40a80f6c207ea06740cd5f4d8f6f0f1ff;
mem[886] = 144'h048c0ef1f904fb06f668fe5ef228f45604eb;
mem[887] = 144'h0ab80c4f079c02cdfe16f042f311f950017b;
mem[888] = 144'h0c350222006fffe8f451f4380732f814074a;
mem[889] = 144'h0bcaf62efeb00c390ced0a75f2e9f30a01a3;
mem[890] = 144'h0f8bf22904ad060afd0d0495fa4effb40d52;
mem[891] = 144'h0e81fa2df719fbf4fb4d06e0f098f67b0731;
mem[892] = 144'hf93e0a8efbedf16d065cfcc10c04037907bb;
mem[893] = 144'h0be5fa920a030ca00b5bf9fb0d63f37af76f;
mem[894] = 144'hf7b804e0f01902810da008c703d707d70256;
mem[895] = 144'hfe050875f9240b58f8e6023ffb0c04be0995;
mem[896] = 144'h0b17f5e6f682fa7efcccfa3508c802d6036b;
mem[897] = 144'h05b802e50751f5ec0a24fbc70e81f514fc45;
mem[898] = 144'hfa2afe61ff5a0376fbb0fd9bf06cf1940f93;
mem[899] = 144'h001d0b0e0dd6f31afcb6009ef9e60d2704d2;
mem[900] = 144'h0cd40b210a88fed307fa0624f0dcfec9fa03;
mem[901] = 144'h09ed04f5fb2c0818fa8cf6b40130ff23051a;
mem[902] = 144'hf3610deb04a0f9f604d50925025c0bfff77c;
mem[903] = 144'h01fe0784083dff4f06e1f65a0f72f7da0de5;
mem[904] = 144'hff3d00ec0a3401fd0b1004550bb4f7a0f7f9;
mem[905] = 144'h06a4f172f31f0c3bf3f1fd150acd0bb3f95c;
mem[906] = 144'h068008ae0343fb56f1f00aa9feccf861f7d0;
mem[907] = 144'h03e9030efe55f217f62ffb41f1f0f05df75b;
mem[908] = 144'hff590903045105c30ab30490f2fcf7d20158;
mem[909] = 144'hf160052b0fc0f1ec0e560bebf61dfb180dec;
mem[910] = 144'hf96b037a044b03be0cbbfa1df5eb00970be0;
mem[911] = 144'hfc7201d404c00439f0d30b840f75f968f119;
mem[912] = 144'hf206ff8b0ee3f7d7ff300981fd5cf3af0433;
mem[913] = 144'h03c30fe40f95ff3909c10ef60c3ff843fe7b;
mem[914] = 144'hf70b0e36f18f040d0372f222f75f04db03e1;
mem[915] = 144'hf7340cb50694fb880486f8e20fa90a1dfb2e;
mem[916] = 144'h0fa30e88fb4504d60f14fdeef20bfb3dfa2f;
mem[917] = 144'h013b0417012e0afaf73700c90e3ef2caf58d;
mem[918] = 144'h07e8fbdefc10efb0003c01770176f1deff3d;
mem[919] = 144'hf13c04fdf6dbf3170340fd2ff696f483ef2b;
mem[920] = 144'hf45c073a058fff05074df0a5f0550e110ede;
mem[921] = 144'hf03efa1bfc34fc00057d0ae4fa4d029bf233;
mem[922] = 144'h0c88feda0ce80c5bfae9001405d3017ef1e5;
mem[923] = 144'h088df967011cfa2002ec0f5c02f2fceffe68;
mem[924] = 144'h015e018dfddaf71d0221fefd0fb3f2b50683;
mem[925] = 144'hfa17ff3b0ed9f1f70ed1f7fff744031d07ba;
mem[926] = 144'h0c54f4ed0241f3ce0f51039b0d02fd000c1f;
mem[927] = 144'h044dfd41f469f125f87af81d040fffdbf1f0;
mem[928] = 144'hf68009b10ef50c1e0f1d0995f258f156f13c;
mem[929] = 144'h07f0fe8af355fa4000b3f56c0534ff660c58;
mem[930] = 144'hf0850514045902770322f480070400f309d4;
mem[931] = 144'h0b5ff7dc01b8f593f1d80d83f7b501f70e98;
mem[932] = 144'h0c4ffd33fb45099005b0f4d7024305a70a51;
mem[933] = 144'h08c0f2bcf254f71205a0f056f724fcb2ff58;
mem[934] = 144'h08760ab9f67ffeea0f01f8dcf893f97bfb8d;
mem[935] = 144'hf1f8015903abf78af5430e6f0caa06aef0e4;
mem[936] = 144'h0153f02e051809ddf60ffcaa071509c6fee0;
mem[937] = 144'hf9faf758f24cfbce0474fddefe91efdd0c75;
mem[938] = 144'h03b8003906a4fe28089c0376083ff4a308dc;
mem[939] = 144'h02f3091c0563f464fb9d05dbf73bf609f673;
mem[940] = 144'hf77cfe3401270987f317fa42fff904b80707;
mem[941] = 144'hfede05540e8c07c4f318060efc75f355f036;
mem[942] = 144'h09af02e6fe58f151fd9b07c70203f8000be8;
mem[943] = 144'hfae6f65400a2f32007d4f95cfdac022efbda;
mem[944] = 144'hfe470bbefe440a1ffbb6fc13f10cf3a107f5;
mem[945] = 144'h0524fa59f9510068f95bf4edf504ffa00265;
mem[946] = 144'hfeb6f30c0b560958f029004ffdc9fe8b0784;
mem[947] = 144'hf443f78df5b705b10eb20290f8acf359006d;
mem[948] = 144'hf78302fbf73df5e6f4f6fc37f53ef830fc56;
mem[949] = 144'hf44f057906df0336f4ddf05cf576feea0224;
mem[950] = 144'h0ae0099b0c87f169fe990aaf0a8b0e0c0a35;
mem[951] = 144'h0c69fab1008ff3dafbf90ef5f6a90a6afc6e;
mem[952] = 144'hf9b0ff1df21f07d50dac03f20d30ef90feb9;
mem[953] = 144'hfb76fd8503cff87d09210edc00720727f229;
mem[954] = 144'hf0aa0b330ddefbcff749febf03b4f90af0b1;
mem[955] = 144'h08220c44f0930970f7870ba20d22fcaaf1bf;
mem[956] = 144'h03a407c40794fd7bf99ef05703d9f3cff35d;
mem[957] = 144'h0721fbf006aa06d1f48b0b78fb5b001807a5;
mem[958] = 144'h0d060b32efea0eaef1240cf5f595fb6f0c2a;
mem[959] = 144'h072bfb7f0579f0db0b7b0cf205e9f7d80abe;
mem[960] = 144'h04f00f02fa2602c109f1f4140bd7f1ef05f0;
mem[961] = 144'hf55508240660f166f05c0c8805830f350cbc;
mem[962] = 144'h0b4508270ea80db4fcdcfb50fd4504650a94;
mem[963] = 144'h06880c1bfba6fd13049c093cf88af12b0309;
mem[964] = 144'hfbbdf2910e86f8dcf55501abf35d05a90436;
mem[965] = 144'hf5df0b7f0955f051fd4b0542fd300a7cfcbe;
mem[966] = 144'hf47b03fe01bff5d7f37d0551fa19f8010730;
mem[967] = 144'hf1ff07a2fc3f011cf2e7f5c305abf13b0e4e;
mem[968] = 144'hf24e07b5fe810a6e0c4e027e0e4b085e005e;
mem[969] = 144'hf905f85b08bc0c9905570636fc26ff5d084b;
mem[970] = 144'h08b4f97e046b0671f25c03d3fb4effab0816;
mem[971] = 144'h065dfdf80de1f65402d1fc330d1f0f4c0ad4;
mem[972] = 144'h0a3709cfff21f807f92f094608f7f242005b;
mem[973] = 144'hf12605c9039801d7f0a4048ef7050db0f64c;
mem[974] = 144'hf977fca8020702be04f0f770f58d0f4f0009;
mem[975] = 144'hf0d90a08fc7401c0f107fad902fdf5340d5a;
mem[976] = 144'h08da0f0100c204660e7505ebf35200ab0836;
mem[977] = 144'h0da0fa6e05e4f794f3160f4c02f7035e05f2;
mem[978] = 144'h0cf6fabe098709180988ff670156f9fdfd56;
mem[979] = 144'hf328fba304d5f4f902f2f16ef2a2f7b3f1ee;
mem[980] = 144'hfbef022cf1c9fbedf5590a3a0ebcf148f901;
mem[981] = 144'h092707fdfebbfc930d8cf773f7df0530079c;
mem[982] = 144'hff16f301f778faf8f0adf3250193f746051a;
mem[983] = 144'h0eedf2660f670537faccfc740f7efa42032e;
mem[984] = 144'h0a78f31707400876f5f5f366f855f37df954;
mem[985] = 144'h039cf15d0eabf0f101b3f7560e81f5caf1d3;
mem[986] = 144'hf0f604d900b3fcea069d0f9d0ad2f3ad060c;
mem[987] = 144'hfc51074806fefbe4f6c50bb9fb31f53cf5e2;
mem[988] = 144'h00eff242033ef834f6e806290662f08f058c;
mem[989] = 144'hf797007e0416026ff6bf0f740918fe56f83c;
mem[990] = 144'h0e8b0b400447fe3606dc0a39fa570caa0c71;
mem[991] = 144'h0dfe06020d43f0ee07110512fea30ce4082c;
mem[992] = 144'hf2720627f495fa81f04e0e20ffe6f73ef0c2;
mem[993] = 144'hf5b0fd6ffa18086c077408d3f664f4e107a2;
mem[994] = 144'h0c93fa9a02710bd4fbcef1d504f5f4560dac;
mem[995] = 144'h0a96f10a007d007af89ffd2efa07f51400b9;
mem[996] = 144'hf1befb93ff77fce70266f811092bfd82ffd5;
mem[997] = 144'hf76df6b1fd48f94e0a44054b063f09d7f8e9;
mem[998] = 144'hf211f91c0a0ffd4dff6bfce8f29bf0d5ff10;
mem[999] = 144'h015ef9e00daf0825086c0e620250003c05b6;
mem[1000] = 144'h0005fa7cf27bf570f8600a3ff4d20d9e0ca7;
mem[1001] = 144'h05b4f341f38901840755f71909c8f6860d5c;
mem[1002] = 144'h0c2cfcbb00e80e0dfed5fdc6f17bf9780e43;
mem[1003] = 144'h016bf923f457ef88facc0622f9940c9a0800;
mem[1004] = 144'hf236f7b7f8b2f100fe8aff3d0f4b0994f70c;
mem[1005] = 144'h05ef017a050ff7d20dcc026b068a06ecf8c5;
mem[1006] = 144'hfa1a01db01410f62f579f918051701ae059d;
mem[1007] = 144'hf064f04c04660298f3cb05a6030608c2fc98;
mem[1008] = 144'h0d64fe4ffaa4021602d00c3504c5f9cdff7c;
mem[1009] = 144'h0dbaf1520426f2e4fd36f4fef094ff1801e8;
mem[1010] = 144'hffae066c0291f43dfe61f5b70e8c0c6503b4;
mem[1011] = 144'h0078f25af394f0cb059e004706ba070ffb84;
mem[1012] = 144'hfa0103d201b5f61906a6fff2f45c0b23fa94;
mem[1013] = 144'hfaa3f38409ad0c30f1c00df00fc5f9d60a6f;
mem[1014] = 144'hf074f143f4430e00ff4fffc403480d7cf919;
mem[1015] = 144'hfefff64905430704ffa8fa38065108e3fcb0;
mem[1016] = 144'hfd7aff4ef2f1f78cff960339efc60af10262;
mem[1017] = 144'h06d50177f8650db9f513fdbd0015f884f872;
mem[1018] = 144'hf880fb3efb38f6a50ca702a0080bf311ff70;
mem[1019] = 144'h0347f33208e9f1f60d2ef77b05d5fd520eb1;
mem[1020] = 144'hf2be000cfa2b096f0c52f410f27cf261f0e0;
mem[1021] = 144'hfa920618fe480cecefe1fa160299f41f0dca;
mem[1022] = 144'hf8240aa7f1b80cb50a1000e1009f00cf0bef;
mem[1023] = 144'hf7aaf7ec00da03a30a7f0c580dd5f6a7febf;
mem[1024] = 144'h0274037f098a0013036a0d4c0e7cf8c4fd37;
mem[1025] = 144'h0cdf0e70026aff28fea2090cff66f0550630;
mem[1026] = 144'h0a21f019f61506b9fb3b0c3ff7ddfac6fa7f;
mem[1027] = 144'hf664056bffadf627045f08dff5690856f370;
mem[1028] = 144'h01e7fe660042fb0d0ead0dc50ec8fb81f0a6;
mem[1029] = 144'hff74f3e0060af6d2003b0fdef7aff3150a0b;
mem[1030] = 144'h06aeff6a0e33fecdfaf205ef0ad6fdfef4fd;
mem[1031] = 144'hf95bf0200ee0043bffc6f517f542f0500de7;
mem[1032] = 144'h0b9ff130f3610b8df90cf2ecfbb7f3d00eab;
mem[1033] = 144'hf86c06840f250d15f07b0a1ff45405aa038a;
mem[1034] = 144'hf26b0687fd34003ff8ebf8bcf06600760069;
mem[1035] = 144'h0be9fcaafd35f875f6f401cef09904b6fd6d;
mem[1036] = 144'h0cfa04ad01a6063d0edcfc220e4702b10256;
mem[1037] = 144'hfdae016df767f5cafb9df041ff900311ffd4;
mem[1038] = 144'h08e206acf460f9bef22b0502fc8105c002f1;
mem[1039] = 144'hfc62f564013c0a72f77bf59d02860eb8f6ee;
mem[1040] = 144'hf1860f300f9e07e10e7e0407f380f157f6a9;
mem[1041] = 144'h0a650dd30863004b0092f372fb76f3e90238;
mem[1042] = 144'hfdfdf8210574fb2a051d0301fe4f09250c67;
mem[1043] = 144'hf3def8e8ff09f09f0c1102e0f7e6f0c9f31c;
mem[1044] = 144'hf7d6f8a3fe33025202c1ff1c0292feeb01c1;
mem[1045] = 144'h020e0070f261f3cd0168fd400100fbd10ae0;
mem[1046] = 144'h0a0af4fe0e7f0e470e630261f0eef4b6f0ce;
mem[1047] = 144'h0de6f7b40dc50c8af9ba0d52fc0dfe48082a;
mem[1048] = 144'h05b206c102bff81505b10bf708ca0ca2fc07;
mem[1049] = 144'hf912fdafef62fb5005e5ff1ffa390717f7c2;
mem[1050] = 144'hfbf709b104ef0466095df2960582fa3fffdd;
mem[1051] = 144'hff5e0344f36c0539fc4306e9081305b8f9a3;
mem[1052] = 144'hfc3004e9050cfc8802c7ffcff64307a7fdb7;
mem[1053] = 144'hf780f1fd0f3efe8bf9b5fd5d0ba902ebfea3;
mem[1054] = 144'hf59300b603a0064cf835f2f5056cff7c0dc1;
mem[1055] = 144'h0e2a019b03a40a7309c1fff9efd0072f049a;
mem[1056] = 144'h0677f2140da6f3aff7c8fa04084dfff9f50d;
mem[1057] = 144'h0e0707400c1f007cffd405f602ad0b340f03;
mem[1058] = 144'hf7dcfff80383015d0f890ad8fbe10c110765;
mem[1059] = 144'h0c68f8c80e8a0ce20652f3e6f64ef8d6084b;
mem[1060] = 144'h0891f84306a90747ffbb0ea6f496fa35fa69;
mem[1061] = 144'h016f0b8603d1f9dc0d400bc8fa780a3a0f7e;
mem[1062] = 144'h09aef7f2004d00eef2ddf39df0b2f87b052b;
mem[1063] = 144'hf049000bf152f39cfb46f114ffe40859fb29;
mem[1064] = 144'h0b88f3e9f4340500f19f0755f7670b28fcb4;
mem[1065] = 144'h0aa509b1f073f429f8fef288fff8ffc9056b;
mem[1066] = 144'hfdbb04c30ba6f99dfc6d0bc603c50d1df7ab;
mem[1067] = 144'hfd98f95ffec3fd5a0dc7faa90c0a062008ed;
mem[1068] = 144'hfa65009c04d30b9d0d5bfee905fc0cc608ad;
mem[1069] = 144'hf6dff4470e7a0a11fc2d0e9ff193fd8b0572;
mem[1070] = 144'hfdc20d2ef690056ef95e007201090696fef8;
mem[1071] = 144'h005ef26101c906ca0a5efcc8f34ef153f7d6;
mem[1072] = 144'hfa9c0f94079b09faf3a0fb20f3a30885f4e1;
mem[1073] = 144'h089200a4f7ce02440db00433f48f053bfaf7;
mem[1074] = 144'h0a3b0ca5034efceb0f63fa8bf6c1f3de0a69;
mem[1075] = 144'hfc2bf6bbf166f1a10268f178fb9c099bf71b;
mem[1076] = 144'hfc3bf23ef70a0d4bfe92058cfda202d5f207;
mem[1077] = 144'hfd20fa4dfdb302b0fdfd024af305f5ed052e;
mem[1078] = 144'hf74ffb8dfc2ffaa0f73af23202390186fe21;
mem[1079] = 144'hfa460deb0d540e630f8df946f5640a710336;
mem[1080] = 144'hfcb708e9f143fb2d0a74f54d00fa02740438;
mem[1081] = 144'hf340ff5f055103a9fa4b04170584ff85f19c;
mem[1082] = 144'h0e590d08095b0086f92ffdebf9a2f3fb0223;
mem[1083] = 144'hfedafeef0c1b0c00f9e0fe6503f70a9ef183;
mem[1084] = 144'hf4a5f1a7f8520500059ff09a0626f15506a2;
mem[1085] = 144'hfdab0d6efb0ff74bf28607b3f132f2cef9a4;
mem[1086] = 144'h085c014e0973f8170d5efe6df452f4c001f1;
mem[1087] = 144'h07f5f33a02d7fb630aef0c9600910eed0281;
mem[1088] = 144'hfaed0da1f31b0329011e02d10f10013c0342;
mem[1089] = 144'hf0f10383fb8502680b990fa80819fbc2fba0;
mem[1090] = 144'hfef0f844f8ccfdc80b99f2d9fa74feaff3a3;
mem[1091] = 144'h04640e1df2fdf9680c44f34309eefeb80718;
mem[1092] = 144'hf19403720aef051ffa2f09acf37d0a7bf8fa;
mem[1093] = 144'hffbe0e090deff44ffe3c09140b0902abf446;
mem[1094] = 144'hf73dfa9c05e2f3bb0be2faaf06e606910925;
mem[1095] = 144'hf412004702a8f88900ba0294fd3d0357f5a5;
mem[1096] = 144'h054bfc65fe6b0b8e0de00705fd96f1200064;
mem[1097] = 144'h0633f2760baaf582f57cfd0ef2151131fff1;
mem[1098] = 144'hf957f67bf6f9fc51f8def4dfff7203de0160;
mem[1099] = 144'h03af030aef26063afb2af4aef45d0f52f08c;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule