`timescale 1ns/1ns

module wt_mem1 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h055205aff793f154f67f040a0ac7fcf5f005;
mem[1] = 144'hf5980ac6f873073b0be50e74f00cf58ff042;
mem[2] = 144'hfeec00bdf05cf462f6e6f02104f1028c01bd;
mem[3] = 144'hfee804b307bc0bdaf1560285f728fdecf3e2;
mem[4] = 144'hf7f6fdedf2c7f29fffa4fac9083a01e2efbc;
mem[5] = 144'hfc6dfe4702c90876042eff92f75bf38efe3b;
mem[6] = 144'heea200d9fc31f820000208f50024f0d5f8cf;
mem[7] = 144'h017bfc2d0a1c0b56ffa30bae099102ac0c13;
mem[8] = 144'hf55a03780bfd0b0f08480c5cf68e0a20fa6b;
mem[9] = 144'h07aa08a2f0f3f6e5078e0c77070bf9a40cbe;
mem[10] = 144'h0a020d77f03bf034f5410379ef2dfde4f0f7;
mem[11] = 144'hf50108ba06b9fe69feb6fa7ef9c9f1c7f1fc;
mem[12] = 144'hfd61f72808c6fe9ff1d5f9fb06370497f120;
mem[13] = 144'h040efb31f2e307e0f52b0631ff4efe8201f8;
mem[14] = 144'hfcea0de50b6f032604d2ee8afc7af01607d0;
mem[15] = 144'hfd2608c5fa26f84103b6f7190d4eefd4fa87;
mem[16] = 144'h0e3d0b0206f406e40e8df5e4fd600c75f638;
mem[17] = 144'h083b0183003807370accef01f0d2f3bef0d3;
mem[18] = 144'h0c17fcf40361033901a90cc80b83f7d0f03d;
mem[19] = 144'hfea0078101d90847f98203bd06410bf90b66;
mem[20] = 144'hf62ef524ff2c02f506ccfa21f532f20503ae;
mem[21] = 144'hf26403bcf810fbdb023c0428fe45f153f779;
mem[22] = 144'hef87f38e096206e3fa400e5a042d03ad0e00;
mem[23] = 144'h0108fb24ff0206e00906f4bc0b9900eafc41;
mem[24] = 144'heee202ad037efb960450f27af5d007e6fc60;
mem[25] = 144'hf9b2031205310341f1c6fd030e04083608ac;
mem[26] = 144'h076701c8fe42092107b6f6fff5fa05bbfa8e;
mem[27] = 144'hf917f7700a210c9af3e2f196ef10ef8af48e;
mem[28] = 144'h0bf2f82bfa100367000a0ae0f08f0b46f27f;
mem[29] = 144'hf53603db0c74f92bffd90c760842f474f9ef;
mem[30] = 144'h083a02f8f955efe10be2f551f24ff4c1eec0;
mem[31] = 144'h0122ff68f4300597f7290e720d9df9400e73;
mem[32] = 144'hef41051b015804bfff8c0851f057f3cdf05d;
mem[33] = 144'h06f00a8ffb97f0630636ff1008dd0a06f7e7;
mem[34] = 144'h06db0addfb3bef6506a507eaf8ddfc6bfa17;
mem[35] = 144'h0aff070af7c0f3300657f644f16af73601d0;
mem[36] = 144'hfbbcfe34fdd3f4d8040a01fd07fc0cde011e;
mem[37] = 144'hfa850d9f02f80ef20b63fd5cf904fe650179;
mem[38] = 144'hf9510dd300d50bc304b4ef700867fa4ffe11;
mem[39] = 144'h0c7c0ad6fd5cf292f20f0b1608e1ff8a001f;
mem[40] = 144'h06000715f85703c1fdf7083507c0f98e053a;
mem[41] = 144'hff9cfe4900db08d7fb290a130bdafa9f0639;
mem[42] = 144'hf11d0b2404dc0875f10efb6a0c9efffbfe20;
mem[43] = 144'hf8da05480458f9b2f21e047df09bef63fe87;
mem[44] = 144'h0cf3ff90fab2f44efe5b0beefc34f004f449;
mem[45] = 144'hfa90f2490a0601e90593f4bbf496f737f4df;
mem[46] = 144'h0bfcf625f0bcf796f0adf26dfe0efc2a0c2f;
mem[47] = 144'h09320131fd73f9ef05840cc2f1dcf908fcaa;
mem[48] = 144'hf4d3f7e3f9ab02b5089ffb670175fd0a0385;
mem[49] = 144'hff0a07eeffc3ffd507ca0b14efde057cfafc;
mem[50] = 144'hffa1fabe0dfaf3210ecdef99f719001c0bd4;
mem[51] = 144'hfa1e04a6f5d104ee0ae2f87e07a3005b02a0;
mem[52] = 144'h02d806e6039cf3f000f00952fb670a24081d;
mem[53] = 144'hf0faf592f156f5f502350418f1c8f99c071c;
mem[54] = 144'hfb2ffbb4fedc07bcf5890bc90123ff1c0b94;
mem[55] = 144'h04acf205f710f9b2072d07e409df0a30f6ae;
mem[56] = 144'hf54af46df4c10ac2f1b70231f6f7047808c0;
mem[57] = 144'h0d93f032fedc0c0f0c8f02c9fcb0fdfcf074;
mem[58] = 144'h08930065050900fcf89405d8fe710a3104a9;
mem[59] = 144'h0761f28df6010839ff16f3bc0666fbe4fa80;
mem[60] = 144'h0d61fc25f444f44a05ed0d1e03920e91fde3;
mem[61] = 144'hf70ff1c3fb43f17dfa61ff98f1d2f1aafabe;
mem[62] = 144'h0d6a0884f87f0255fa6b08f8f3ff0d610db3;
mem[63] = 144'hfc47048c040bf2740c2d0b7806d6002804f1;
mem[64] = 144'hf3c4f56def95f0b1f982fbe1094d01ae0675;
mem[65] = 144'h0de007ae07dcf6b9f39204b00842f44e0294;
mem[66] = 144'h037af236f5dbf7bcef9e02b4f50c0aa100d9;
mem[67] = 144'h08eef3110eb6f979f361f9ce0359fea8f674;
mem[68] = 144'h056808faf1fffd00f42105420c1cfd9e0f98;
mem[69] = 144'h09280e31f208f278f443f99f0c5ffcef068a;
mem[70] = 144'hff1f06610856067407e5fa3708cb0e35f555;
mem[71] = 144'hf7fefadb0536075bf3b500890414086b080c;
mem[72] = 144'hf4d0031df2b0fc8104180df806740dfdf1e0;
mem[73] = 144'hf63bf0fff796023a060f0986fe01f59af091;
mem[74] = 144'h0f250a97f6c2f78b00eafb0bf9ac08ab0891;
mem[75] = 144'hff1afb30fb33046007e80438036908650537;
mem[76] = 144'h02e5f3e3ffce0be3ff90f3c50c5f0b73f2e0;
mem[77] = 144'h0e19f657013f080a0d7700d902cef1310756;
mem[78] = 144'h0b1d0c26fd84f3f9fe3ff9d2f1510e180a34;
mem[79] = 144'hfb8df6b2058c0eae0322036ef1680c1d09e2;
mem[80] = 144'hfb98f52d04d3f769f563f27efd1bf515fde9;
mem[81] = 144'hf7f207bbff85077f0e8bff90ffbc0252f10e;
mem[82] = 144'h0731f2edf1aa09d607a5f1b1f880fe60fcc8;
mem[83] = 144'hf731004104110361f17f0149ff74f81df87a;
mem[84] = 144'hf180f0a70768f5caf063f2f8043afeaa05f9;
mem[85] = 144'hfc32fc2a0419f1b30b39fbc5f13408daf106;
mem[86] = 144'h02aa0699fa6c02ac06570a76fe6004bf061b;
mem[87] = 144'hfd01fe920ab703de032ffc00feaffad3fcea;
mem[88] = 144'hf6faf03a068308a5f1c201970b9df7b80366;
mem[89] = 144'hf81a05b8fb1bfceb09b5f7cd0227fff7f6c1;
mem[90] = 144'h03250e19f257fb1a0085fe320779f5a1fb5c;
mem[91] = 144'hf5f70e8bf40e05def5ca0e08f2d7f179fa82;
mem[92] = 144'h07a2fe09efff09650843f40b0d45f691f74c;
mem[93] = 144'h03b2ff7204290370fdbdf478efeef191f579;
mem[94] = 144'hf1b1059bfb2d0d19081e0e89f21af3090534;
mem[95] = 144'hf931fb37f93a026ef8bbfe2af3250194f5f3;
mem[96] = 144'hf40a032ffda70d29018805670e2608dcfbd8;
mem[97] = 144'hf1cc055c0b88f5b2fa2203b60981f084fbb8;
mem[98] = 144'h0f77f28603050a6f0f080b240fb2f1ce01f2;
mem[99] = 144'hf73d024b0bf3f7bdfb2cf007fa3f0167f8dd;
mem[100] = 144'h072efcdcf77a00920cb40ea1fe760a3f0a3f;
mem[101] = 144'hefeb088904390b10f8e0f7a7f2a00c0505ee;
mem[102] = 144'h05caf6ce02a4fecff4fc00890258007f024b;
mem[103] = 144'hfaac0507fd6dfaad03caf2d0f5be0a840e3d;
mem[104] = 144'hf2c7f189023d050b0ba9ffa7f52bf089088f;
mem[105] = 144'hf6a6f24702750b44fcb404460c8ef078034b;
mem[106] = 144'h030df5960b2a0317f2edfa71fd440ee602dd;
mem[107] = 144'hfb19021e056f0c5e04260fbbf4720d550508;
mem[108] = 144'h04c50240fa7cf28e0738f7470cee065bf93c;
mem[109] = 144'hf323f4a4f6b5013d033f0d07fc66fcb205b9;
mem[110] = 144'hf244f37a028806c20659f5d20b15fbc10d39;
mem[111] = 144'hf6a30b7dff5c05b3fe6407ebf461f6f60c46;
mem[112] = 144'hfae202a1f539fa4cf5c4041101a1f8810d5e;
mem[113] = 144'h0cd0fd98fa45fdeef057f8b30895fa0a07ee;
mem[114] = 144'h091405510419f4f9fab00f8f09d50b5a0d75;
mem[115] = 144'h0725fd0af7ee047102b1fb46098ff47608c3;
mem[116] = 144'h02cf06b1f5c30b4ff5990c9e0ab500800be9;
mem[117] = 144'hf8ddfbbc03e90a7ef651ff63f6e7f6f1f873;
mem[118] = 144'hffc5f76f022801fdfdde0a480b5fffb109e4;
mem[119] = 144'h0425f0dd0975f089fe69ff63f2b40604fa07;
mem[120] = 144'hf07e08e0f80b0be5f9fff140f8adf1d80185;
mem[121] = 144'h07f7f0870e5b04d20699f3550059f2c20659;
mem[122] = 144'hfddcf945fc3a070d0a31f408f58bf57af066;
mem[123] = 144'hfa1af3ef0455fdc301a10dea01b30be9008f;
mem[124] = 144'h0e09fb9c0861fbccfc40fd440c8f039603fb;
mem[125] = 144'hf69df072f6d5fa5c05350355f7a4043bf9c9;
mem[126] = 144'h096e05aafa98fceff9cefc1d0a60f7d4fbdf;
mem[127] = 144'hfccdfa0cf7d0f5730ad5f849f17d06dcf657;
mem[128] = 144'hf966027b0f99f77d0017fb780569069b0729;
mem[129] = 144'h09880387f279ff530a1dfdf2fd7ef212f562;
mem[130] = 144'h0552fa68fcfc080ef4b9f9d9f1a5f8b3f8a4;
mem[131] = 144'hf844f8f0040a0e0c07f4f2020270f1c70967;
mem[132] = 144'hf578fd26f2e3f64cfc3c031af4120f01036d;
mem[133] = 144'hf14cfa8a0107f94df2f5f949037e0c2207e6;
mem[134] = 144'hf192f6ce0c59f06d065d04200b1e0d400fe6;
mem[135] = 144'hfe140fe7072ffd9b01a3fb26f2270eac09a3;
mem[136] = 144'h012ff85704e900eb045cfda8f7f303250cd8;
mem[137] = 144'h0b1b0efc0a79f65e0a21ff1af89c04c7ff78;
mem[138] = 144'hf60e0ed7f7280769f94c02730d6c0eeb0253;
mem[139] = 144'h038efa90067ff80dfd34f3430f3506590a37;
mem[140] = 144'hf179f9b006f0066409c9f573fa0af2a70e8f;
mem[141] = 144'hf84af196fa86f8ec08eff64ef39ef1b5f12f;
mem[142] = 144'h09f80b56f5e8f17509c1024dfc8b09acfd8d;
mem[143] = 144'hf65aff51fe5b0f48fab302ec0786f703fe0d;
mem[144] = 144'hf2fb078ff81cf36d054efc41f2da074bf530;
mem[145] = 144'hf006f4cd08cc050c0e920376f4370a1afeae;
mem[146] = 144'hf938f1def936fa2503790278f7270998ff64;
mem[147] = 144'hf1bafa60f6f6010efcb1f8d2083605c60ea8;
mem[148] = 144'hf98df50ff2b0ffa8f14d07e90333f342ff22;
mem[149] = 144'hf8fb0709f2f10bfc037308020ac50acf076d;
mem[150] = 144'hf91e02310636f5720a1bf6d800050a99010a;
mem[151] = 144'h0084005c07a30da2f7df0913009e007afbb7;
mem[152] = 144'h00400cd3052c0979f4300a00f5fcf51affc7;
mem[153] = 144'h0662094a0b9206410aaef5fcfc21f57903bd;
mem[154] = 144'h073a08abf8d000df0e9d0b28079f029c0a5b;
mem[155] = 144'h0de1f1830b2c00f0003001ce084ffaf4fe8f;
mem[156] = 144'h0e3bf1dafd31f0b3f442f0b5067df3fff59c;
mem[157] = 144'hfdd70215043df0e7f702f8d8fa61084f09d6;
mem[158] = 144'hf481fd6b077307f1eff5f9f900a7f0800a71;
mem[159] = 144'hf30808200b60054907e3098ef4c000ba040c;
mem[160] = 144'h012af3b9fdf90aa60e93f3ce0c7d015af937;
mem[161] = 144'hf5ef057b0cfa0ad0f42bfc20023b06e00372;
mem[162] = 144'hfc27feaf001404d6f48ff2c009d40aa2fef8;
mem[163] = 144'h0693f2b1f5b40966fd7af71bfd0efa79079e;
mem[164] = 144'hfceaf7d306e80bccf7f9f8ed0c9906e6f81d;
mem[165] = 144'hf35101ec0d2a087dfd64f4c0fc940845fcbb;
mem[166] = 144'h0c2c05e101c6fd9bfb42f498f23afe7ef59c;
mem[167] = 144'hfab005940c780dd50f17fa4405830e040fbf;
mem[168] = 144'h0a6d08b2f6b2f6eaf13df8810dcbf297f91e;
mem[169] = 144'h0501f1be06d800d2ff06f89109350afe07e6;
mem[170] = 144'hf19f0d8901cafd72074af98df159fd5b0591;
mem[171] = 144'h0ea3f77af1edfb66f1f4fe91f7abeff9f5bc;
mem[172] = 144'hf1e80b87ff3df512fe5bf0c90e93fbe40cc5;
mem[173] = 144'h06a6f7a80b52f96c06d2feaf01a1ff4bf69e;
mem[174] = 144'hf88e0a90f3480076fa310835fe3ff2f3f1e4;
mem[175] = 144'h04a6060bf0a1fc27fc61ff48009b07b8f1d8;
mem[176] = 144'h068dff62f3d90305f06002aa0f4e02970293;
mem[177] = 144'hf41005440d6703120b4f0caef761ff97f183;
mem[178] = 144'hf3f1ff660b06095a0a3d0ac8f7cbfb2a069f;
mem[179] = 144'h09ad07c1ffccfb8dfea107b4f90b053e0f0f;
mem[180] = 144'h04630540024008cf084ef803fc84f00dfce1;
mem[181] = 144'hf568fe70fe7f0bfc055af36e0200f33e0b66;
mem[182] = 144'hfa1f019b0e36ff8af0e9efcd07e1f074fadd;
mem[183] = 144'h0587fe02f170fc170efaf05eee9a01ae0cd5;
mem[184] = 144'h06cffd8f01600b35f3330052f279016705c3;
mem[185] = 144'hfec3fc750f1d0c000c45f1a2009df68df9ac;
mem[186] = 144'h061bf437002afea703690b4f0830fb7e0996;
mem[187] = 144'hfeb2037df9020e00f21a0dd701c1f78a047a;
mem[188] = 144'h09ab0158f57af4330092fd5af67b07f7f59f;
mem[189] = 144'hf584fc090803fc760f0f0afb0e67fc6e0a4c;
mem[190] = 144'hf9b00df3f1b9fa81fe060a160d53090ff47d;
mem[191] = 144'hfcc9fed4f523f55ef81df41bf25e0b4bf57d;
mem[192] = 144'h094408010190f5e5f5b408b9027af5bb0667;
mem[193] = 144'h070a0b07f8c10de4f1ef0ec0064bf514fd78;
mem[194] = 144'hf95f0cda03a5006ef630fa43ff5af0f504ed;
mem[195] = 144'h0f91f7e0056cfdcafd29fd11f836f0420541;
mem[196] = 144'h014003b2fb340b78f711f7a0f0710edb0817;
mem[197] = 144'hf93ff3f80f2af66b055d0924022fff7504a0;
mem[198] = 144'hf6ccf3040c6af1a9fde70e7d0e400e59f6d1;
mem[199] = 144'h0179f5e6fa1f02a40e92f9d8f7b30f820ea5;
mem[200] = 144'hffb50d810000f31afa82f62aefe908bbf608;
mem[201] = 144'hfff003a90a88f7e7067af158f3d209adf441;
mem[202] = 144'h04df09b4fabf05fc0d01fbfc027cf43bfd24;
mem[203] = 144'h06050cbdfbb70a0709b507290b0e0c07ff0d;
mem[204] = 144'h00edf1230b93f27ffbeb0897f2b90170051d;
mem[205] = 144'h0f5bf25ef9070932ff30f830f1b30153f9f7;
mem[206] = 144'hf21a02f701d2fc44f6d5029ff773f160f09c;
mem[207] = 144'h0b74f4f2f0d50fbbfa110707023e05e40bc1;
mem[208] = 144'hfc60fdb90df7f61e02430362f23c0c6e0144;
mem[209] = 144'hf450f9300a5c0b270ec5f51cf3cd014d0243;
mem[210] = 144'hfd3e0f15f11b06d5021c05e3f5320eb7feb9;
mem[211] = 144'hfae3f53a08e8fcf20cbff82e09aa05c60399;
mem[212] = 144'h0be4fdd4031800430ceef55f0205f1270162;
mem[213] = 144'hfb18f9160e8cfbdcfab1f51bfccff650fce7;
mem[214] = 144'heff5f4a203a8093bffddf2c8efeafd5f0e97;
mem[215] = 144'h06f500e1f87f0b4b0b1b0849067e094ff1f3;
mem[216] = 144'hf5070768022bf546fad2f043f7d0f95c0aa4;
mem[217] = 144'h01f202e9012bfa0e077d082d066e03c606df;
mem[218] = 144'h0b5a032a0081089a0609f893fcfef738f31f;
mem[219] = 144'h0ab4fd6801c10e1df8ebfc970cd5f764fb6d;
mem[220] = 144'hf396f87bf0d9fc19f90902adf567090d0485;
mem[221] = 144'hf636f7ebf5350f03f858fa6ff78e0d11ffc6;
mem[222] = 144'hf36c05630c34f0dcf73201f5f827fc72002e;
mem[223] = 144'hf07a09b0faf8059ef71ffd13f276fe4afc48;
mem[224] = 144'hf59bf8b5facf064a05f00e50fec800adf2fc;
mem[225] = 144'h0ad905c3098f0c0f025a004b03b30c21fc37;
mem[226] = 144'h0587f117ffb807670a0c0c5bf28cfc93f3b3;
mem[227] = 144'hf65501480b79fbfcf18bf50bf978f697fd5f;
mem[228] = 144'hfd4b0350009ef94e04280770028cf559f984;
mem[229] = 144'hef7df5e8052df9990cbbffa7fecf0572ff2e;
mem[230] = 144'h00ac0deb07eff9880a46f7cbf20305f90c26;
mem[231] = 144'hf2c4f4f50a7b0a22001bff8a0643080afd12;
mem[232] = 144'hf1350c69f7dd0013f0ea084af6090a370739;
mem[233] = 144'hf001faa5fa990738ff0307affb2c05cbfe4e;
mem[234] = 144'h0b0701620d5ffdbf0c45f03afdb2f74b0ebc;
mem[235] = 144'h0e92f18a00c2f0edf03df70f043b0316f545;
mem[236] = 144'h093df8cdf7fe04e20eb507a0f89301c90dc7;
mem[237] = 144'h0d3e0633fd55019ffa62f5f3076705ee0ce8;
mem[238] = 144'h0c2bfa030aea086903fafb29fee7f09a0570;
mem[239] = 144'hf3ae04b9fe5902b5f639f11ff432f69a0c37;
mem[240] = 144'h0803f9e50cf10f1afafb0b84f70f0f4fffd7;
mem[241] = 144'hf3d00ea807ce0f9e08d403ab02a6efb3f865;
mem[242] = 144'h08d70c30ff050d5003740426f52400d90144;
mem[243] = 144'hf665029cfe63fe1f0189f9f0f5e80d270515;
mem[244] = 144'h0dbcfe0e0d6cfe63faacfde7f2e30386fde1;
mem[245] = 144'hf9e4041d0ee5ffd70c780ab208c7f79df022;
mem[246] = 144'h0fe2077f0b04f2b0fb90f9670170f87b0d76;
mem[247] = 144'h04e708d3f508f96e05160a8a05130df7f75d;
mem[248] = 144'hf1470db2f90c0059f6d60f160cb008cff49e;
mem[249] = 144'hfb190f08f5caf86e0ec8f28cf5730e91051a;
mem[250] = 144'hf825fe24fe7af13706a90d41fc010f77fd19;
mem[251] = 144'hffca0a8c0c49080df452042603940e35039c;
mem[252] = 144'hf8bd02caf7a10222fdaff18ef6fe0111fb2c;
mem[253] = 144'h050600daf54dfd56f5e405a1f77a0f15024d;
mem[254] = 144'h069909f70a10045302f20ed30371fdfcf34b;
mem[255] = 144'hf1930eee06f0fd960571006603f4f6e2f9ff;
mem[256] = 144'h037a0b4cf7f30c5dfa840de8fdeafd490f1a;
mem[257] = 144'h0418f89e0d34006801e6f06b0985f4410890;
mem[258] = 144'hf8920c21fb990cdefe25f6ea0e9ff430fc1f;
mem[259] = 144'hf48d05fef48efc85fa2a06d6041d0d5afcb4;
mem[260] = 144'hf3580dd5018b0c8fefb8f2aeffd6f6c8ff3b;
mem[261] = 144'hf527f59bfae20c0e0c99fb3907b0f94309d5;
mem[262] = 144'hf1adf766f4ce03be07cc03c303b7fe04f00f;
mem[263] = 144'h06b7f20e08e50fbf0d51f453f228f9e6f6f9;
mem[264] = 144'h0b59fa6ef8290aa7f13d0441fbb3fea6f140;
mem[265] = 144'h0bd0fb6cf0cd08d40ed3f895fcadf1920c5b;
mem[266] = 144'h0767f719f1d0f3a7020ffbf1f88f039d057b;
mem[267] = 144'hfddbf0faf750f8a2fbe602b20914f03f0c63;
mem[268] = 144'h02dfff4c0f39068ff6bd013aef67f5fb0ac4;
mem[269] = 144'hf996f457efc40c7ff809f35ef9dd05ea0839;
mem[270] = 144'h0ba703f6ff7709e9f01b054dfbb9f72d0ee5;
mem[271] = 144'hfbccfb8b0a5f035906a8042cf4d2038b044d;
mem[272] = 144'hfb5dfe740289fd92ff7d0c3e08e20338f1e7;
mem[273] = 144'h0ee1fcfef5a40869f7d0029a09ddf6b1f789;
mem[274] = 144'hef56083b0e8a0ddaf1c505c307ac08b3ff91;
mem[275] = 144'hf3fef9d203b803fcf8950d2f0445f61f07b4;
mem[276] = 144'h04840308f5760401fb9cefbdfe82fdac095e;
mem[277] = 144'hfbfb0d11fc60ffeb0a63fb8f0d65f9680558;
mem[278] = 144'hf747ff4f0367f193fab2f94eff8d04b8f437;
mem[279] = 144'hf54d011ff124fa6af78bf8c0efc2f06aefcb;
mem[280] = 144'h05d10e6befd80ec00f2f0daf0b94fb7bf049;
mem[281] = 144'hf352030704bff65e0ad4035af8da07e7fdef;
mem[282] = 144'hf4b5f7d4011bf4edf3510b2ff1090770fc9b;
mem[283] = 144'hf669fbe4fb52f68a024a03840996f434f01d;
mem[284] = 144'h0608f8c60b02fd6cf7b4f8e30729ff2c04a4;
mem[285] = 144'hfb7400fc07f2fdebff390dc306cdf90bf93d;
mem[286] = 144'hfa85fd31f224f41beff005fb07cb0c8e049a;
mem[287] = 144'h0e75f3240e670eb6089a0acef9840ddcf96b;
mem[288] = 144'hf6e6f181f4a101240ecff50af8c20e99f8d9;
mem[289] = 144'hf3f60457fa6bf8faf9a20681fa36f4b6f627;
mem[290] = 144'hfa7ffe2b09f20d30f7af0569fe350188f160;
mem[291] = 144'hf3ae0776f024002304f5096d0952f736fc57;
mem[292] = 144'hf0360dd6f3e0f7cd04020a100094ffacf9f7;
mem[293] = 144'hf276f8a2fcfc01f502e4fd1efbae0d440ae3;
mem[294] = 144'h0436f9c50c94ff6ff5fa088f0bacf4d8f79d;
mem[295] = 144'hf720f84f0203f75a0d9307d90b35f7140c2e;
mem[296] = 144'hefa80703077009550927fc8a0799f0700286;
mem[297] = 144'hf12af07c0d20f30f0ef402a5020f09f40e01;
mem[298] = 144'h0d12f9c7f21a0aa4f8d1f432ffd6079cf414;
mem[299] = 144'hff4507b70f5dfffa0fecfba70da4f7d203e3;
mem[300] = 144'hf107f81a08580d290bbc003a0efaf4060e05;
mem[301] = 144'h0392f2fcf26c0560f24c04ef00bf0d00ef72;
mem[302] = 144'hf93600740e5a02acef58f7eff30dfe43043e;
mem[303] = 144'hfd0d00bcfa9ff09c09b40f140e7000bbfc00;
mem[304] = 144'hf1920135f41409b2063af21ef914030afd3f;
mem[305] = 144'h01c1fafa0b1b0251fa9707ecff12f2e1f0c2;
mem[306] = 144'hfccef1760b90f91f082008c0efe20924021c;
mem[307] = 144'hfb36f795fc35f882fa59facd099d03f3fd98;
mem[308] = 144'h02b5f20209a807e50dfdf088fb2705950c86;
mem[309] = 144'h0b1e085405e3043ef3dd0e0a093d0bcc0346;
mem[310] = 144'h004803bbfc5107aa09fbff77fbab0ae0f55c;
mem[311] = 144'hfadc09aefa24f0ee066ef0baf84006d60213;
mem[312] = 144'hff2b0b14fed6fbe6f6a50edc03b005defcc6;
mem[313] = 144'h0c4801180209fc610d8a082cf1a2025601b1;
mem[314] = 144'hf32f0aa405ecf4cb0b67067d0919005ffd5e;
mem[315] = 144'h08def227f836f1faf474fea3074805dff877;
mem[316] = 144'hf6d000360d2800acf335f7960a23f4090348;
mem[317] = 144'hf9c1f33908d0f08dffd2fedefa8bf5e3f06a;
mem[318] = 144'h05d9fd0c0532f252fbf9fb55feeafe47f7d1;
mem[319] = 144'hf28b08ae076df35707620212f2da0ce4fe0e;
mem[320] = 144'hf660006ffa720099f13508e30d49f1f00ef2;
mem[321] = 144'h093efdb703f7ff9a0e64fb4b05dd0763f5ba;
mem[322] = 144'h0f34063cfee8f3dc0437facaf389fe3cfd6a;
mem[323] = 144'hf996f7cd0505f8830ea604380ced0ca6f4b7;
mem[324] = 144'h0acf0c4202b7f8d50a63f7e20670f9e1045e;
mem[325] = 144'h0e4a0ca2f2f5f9c80a150f4bf5400879015f;
mem[326] = 144'hf003fc6ef9aff2c20ac6054f0ea4f70cfa0c;
mem[327] = 144'hf16b02da0cf3061809c30186f44bfb9f005a;
mem[328] = 144'hfa3bf1ca09adff1af518f61a01870b40fc30;
mem[329] = 144'h0b620a8b05c3ef99f649fd5ef69e07cd02bf;
mem[330] = 144'hf7da0e9f0846f8d20b69051af0ef09a60247;
mem[331] = 144'h0e13fe19fa450526f02803170f59f22d0f65;
mem[332] = 144'hfe82f0ef0404ff6bfa5e03d807a20c2c00d5;
mem[333] = 144'hff19f0d70d660095073f098b028a096ef477;
mem[334] = 144'h01ff0baa045303d907330e9af7ad0377fecb;
mem[335] = 144'hf212f9edf1250c56064905a00f5206520139;
mem[336] = 144'h016ff269054e09c0029802210218f9fbf2ad;
mem[337] = 144'h06950475f6f707c902ef001af4790dbdfa12;
mem[338] = 144'h0d42f05208a70895fdbafb00f54efe69f427;
mem[339] = 144'hfb850004f15107a9005f0df7f6560e3ef492;
mem[340] = 144'hf626f05df965085d07d8fb14fc41fbe0f302;
mem[341] = 144'hf4fbf3e8fc4d04f4f3f5f055ff86f1b9fe9e;
mem[342] = 144'hf1b5f1140989ff67f444057af649fa54f6fa;
mem[343] = 144'h02a5fa1901b30711efc6fdd4041df520fe7f;
mem[344] = 144'hf5a109e2f8570af9f450f0e203f8ff09fcc3;
mem[345] = 144'hf1baf10b01e205b5ff9bf712fd47f6750fe3;
mem[346] = 144'hf3060130f610f1230647f35dfc4202a3f2b2;
mem[347] = 144'hfafaf2740bfd09adf238fb85fd42f4e40898;
mem[348] = 144'h08900d040ab3f36a0bbaf4ae0f4d0f35fdc1;
mem[349] = 144'hf769f8cafae9ff2bf49f016cf653fa240781;
mem[350] = 144'hfa0bfa5c0f37f277f178f29ff70306cef198;
mem[351] = 144'h073f075efd4301690e6ef512ff83f2e909e2;
mem[352] = 144'h0d5e0677fc78051e045ffc110198f7590e67;
mem[353] = 144'hf62d0795faf8fe41025bf17e06270e480013;
mem[354] = 144'h0744090c06ef020f0d0df3acf6b4009cf26c;
mem[355] = 144'hfa35fb0f0be905780c1b0636f49f0ea60514;
mem[356] = 144'h0b27f6d300c3015efd8601850961fe6b046c;
mem[357] = 144'h03730da3f687f9adefb607350b07f4b20ae6;
mem[358] = 144'hf951f656fee00467fa2307e5f41bfd43fc0d;
mem[359] = 144'hf6fcfa7a029b078afc33f5e3efb6ff4f0f8f;
mem[360] = 144'h0dae0eecf4740d4806c1f833fb120661f873;
mem[361] = 144'hf4cdfd2b080a062e00cc0b3af84ef00b0d43;
mem[362] = 144'h008f0ddc088eefe6048ef0120e7af392f8eb;
mem[363] = 144'hf59fff82f551000efe4f09000303001c0b7d;
mem[364] = 144'h081afbc0011e0187f73305c4f81bf55bf7e3;
mem[365] = 144'hf4ab0b5708e4ff3ef759fe0808f7f990f02e;
mem[366] = 144'hfb06efff01e50d9201c1f0500b5cf39df78b;
mem[367] = 144'h03eff6c0f1990f27fb2602e6fe3d0ee90d13;
mem[368] = 144'h0dd402f40be60cdf0f260de30ad1f58e06ab;
mem[369] = 144'hf27ff584fd37ef500b1202a70f13fbfaf24c;
mem[370] = 144'h09b7fdff07fcf028f1caf3aff1810e29fac0;
mem[371] = 144'hfbb8f31df4700d1d005b079205eff5def448;
mem[372] = 144'hff5a0f8103670dee0a1afe53ffb9f95bf457;
mem[373] = 144'h0d57f7650edd044d03b3fc55f543050801bc;
mem[374] = 144'h0c18f8dcf5b50f9b055cf811efdc07ce0f7c;
mem[375] = 144'hff98f4370869f32af1cf099c0031f228f09c;
mem[376] = 144'hf1fc02c5f27df623fda5f3abf2f8f5ec010c;
mem[377] = 144'hfc52f5dd0ad5f3dc08ff0775f4c5fbd6fae7;
mem[378] = 144'hf792fab60ca8ff1df848f96f0b7f02bd0ee7;
mem[379] = 144'hf3c401c8061eff65fb25fc3309f5f71afe41;
mem[380] = 144'hfb7af32c01a2f39cfbaf08cffef30832048f;
mem[381] = 144'hfe710cc207f602b8f592f391f1d9f607fb3b;
mem[382] = 144'h049f071a0618074b07eaf94cf3a4fb8e0bcb;
mem[383] = 144'hfa9eff4b0ed203e20de10a83ff4d02f5fa62;
mem[384] = 144'hf73cfb770832f1de028cf5e403c80d6505e4;
mem[385] = 144'hfc4c0a08fdd4024703d407440962f9660d90;
mem[386] = 144'hff20f167f3d505bff38b09bcf20e094d0e9e;
mem[387] = 144'h05e70dd80a17feca0f350206078bf5d60e09;
mem[388] = 144'hf745f5c204d2f991efb706ba07bdf4b4f7b0;
mem[389] = 144'hf0b006970a70069c0df309f00684038ffe87;
mem[390] = 144'hfe2afffb0689f4ad00bbfccb0a15fe7bf53d;
mem[391] = 144'hf55203b0f4fef18b02e9f12a0b39f10bf083;
mem[392] = 144'h0ee8020c08170e7f0c7b00e0fd38fb5afe87;
mem[393] = 144'h09c90060055efb25034208f5f15b00ec0420;
mem[394] = 144'h00950671fd97099ff383f9710cd3f428f8ab;
mem[395] = 144'hf8f1fd2505740f3ef32bf049f1d0f9c4fcbe;
mem[396] = 144'hf6f0fc02f19cf759f4c0009af8c8efc8fd3c;
mem[397] = 144'h0bd4f6f1fd0efc310a670ed6ff92f1270d59;
mem[398] = 144'h029c0db90174f34100d6f70df4030fb2f51b;
mem[399] = 144'hfb2306fdf3b60e42f8ba026dfb3f071a0db9;
mem[400] = 144'h016d0cf30f82f186fe6df3f201f5fe1e0ec1;
mem[401] = 144'hfae507bf0ae208630e600eb60efffa17f672;
mem[402] = 144'h0ab6f660feb1f7590af501c605acf7c0f21e;
mem[403] = 144'hfa0803740d810f9f073ff8b1091e0a230d30;
mem[404] = 144'h0691050809d2fee6fc870619f7acfdad029c;
mem[405] = 144'h0b16f507fdb6f36104050241f82a0aa105d5;
mem[406] = 144'h0af30284fb5df6ad0d270b530bf4f13bfc38;
mem[407] = 144'hfde8fefcfb8ef06afd5d0c400486f3680201;
mem[408] = 144'h04760278f297fd2bf119f0f1f29c0ebaf2da;
mem[409] = 144'h086c078b03a0f4c0073d08b9fac0fb930790;
mem[410] = 144'hf36af032fd170c310973f369f85ef51d0ac8;
mem[411] = 144'hffc60279f3f10bdbf085096a0793f535fb71;
mem[412] = 144'h09bf0658f2640c30f498010505500553089e;
mem[413] = 144'h0f9a0d8701a404b8f10b099bf750f29b05fd;
mem[414] = 144'h0e99f8a70c8efb47fd2f0d040736012b0019;
mem[415] = 144'h029c04b2f390f5c7f57a0e1cf0a90a11fe22;
mem[416] = 144'h0750f54cf117f727f88c09bffccaf9a305ca;
mem[417] = 144'hf6b2f7e8fc140b5bf7810ea50a80fddb0c5f;
mem[418] = 144'h058df835fbd60a73f3f30ec40151044302c5;
mem[419] = 144'hfed7ff1ef7ed0caef002fd1b0009001f066b;
mem[420] = 144'h02070c5f0c4403f0f5f303d7fd62eff303c6;
mem[421] = 144'h01bf0b61f31e0ea70bbd0a47f3aa0ecaf28f;
mem[422] = 144'h02ed09b003e8f9eefc78009cf7f9fd1501ce;
mem[423] = 144'hf78bf687f6be095b00bdf1fa0088fcb9002f;
mem[424] = 144'h02a305fcf9cc0a37f957073cf701f3ec0650;
mem[425] = 144'hf63c01eafa72f449f32ff7990156fd540c36;
mem[426] = 144'h070d0055f183f38002c6f74cf72002aff7ba;
mem[427] = 144'hfa8efe61f43ef17af2d10b69f5760cba0f17;
mem[428] = 144'h02e3091efc870c48fd16f536f2daf90f046b;
mem[429] = 144'hf3fe04aafcc5f1610e8109bcfe5b0669fd49;
mem[430] = 144'hf3cdf03e05b108f007480185f5dbfe76f0dc;
mem[431] = 144'h0ee0f01e0061f684f1c4f54305b0079dfc33;
mem[432] = 144'hf7c90df0f583fa180253f9960e4809f9f5bc;
mem[433] = 144'h0e75f2a403e0091d006e08aa03b5fb0ff9f5;
mem[434] = 144'hf933feb50dcbf78d0c6c0919f92cfeeaf680;
mem[435] = 144'h008d0b8af0bff3e30ddff05b0cc40deaf04b;
mem[436] = 144'hfeb0f2dc009b00d1f15cfe68f98df111fc71;
mem[437] = 144'h0452f26ff2ac0afafbeff3880beefdab0d3f;
mem[438] = 144'hf3ae0f1afcd7f30dfd5402fa0871f145f3b6;
mem[439] = 144'h0d27f7f1f53af67b0bef0aa502cc040af8c8;
mem[440] = 144'h0a010ae20ceff01b0787f8dcff69f0d80534;
mem[441] = 144'h0d53f10af8f1f21efe17efc10a88f3240f02;
mem[442] = 144'hf5ee0ecf0741fbb2048ffa65019d0a42f43e;
mem[443] = 144'hfe20fe21f0580dd7057408fbfb1609abf797;
mem[444] = 144'hf89af3f10b99f132ff92ff61085ffe86f0e9;
mem[445] = 144'hf85a0e9dfae500c60c3a0565059408a7f695;
mem[446] = 144'hf9b3fe06f7e20efff598f0b3f2a80ca1f3eb;
mem[447] = 144'hf079fa040534056e0d56f8040982fb1d0b6f;
mem[448] = 144'h04b7eeb60967f3670d91f215f7a40d6408d2;
mem[449] = 144'hf900f8990148f4e50a52fd20f34504f00853;
mem[450] = 144'h0a27fc750e6ef85603abf490f753ff29f3cb;
mem[451] = 144'hf704f8b209370790fee1f037f30b0d02f3c6;
mem[452] = 144'hfafbfa3e098f0a2d0517fd11f5e1f8faf3bd;
mem[453] = 144'hfb2701400cb406f604abf91c0132090af726;
mem[454] = 144'h0312fe62f266f452f2a701f709d6f08aef7b;
mem[455] = 144'hf990024b0eb7f5fef330f5ab083f05c2fee5;
mem[456] = 144'h0a35f73b0577f316f727fd5ff97cf05cfdfd;
mem[457] = 144'hf44f0c090367085ff6f80a48064602170617;
mem[458] = 144'hfbd3fcaf0c9e0f5efbfef670fad5fc750f08;
mem[459] = 144'hfaccf8740448fa7f0919f8c20307089ff54c;
mem[460] = 144'hefa7fa00ff2d02600a9df4c1035ff3b7fd4e;
mem[461] = 144'h0652044cf1c0f6520e29fd1309ccfcc8f311;
mem[462] = 144'h06bb0e720a1df333f4810ea8efa1f868efd3;
mem[463] = 144'h05ee09d30f7f0efd003d0b340cff0b01047e;
mem[464] = 144'hfb3f0d2e063ff48f0d7909e4054fffd90701;
mem[465] = 144'h0772053b094407f90f08054af21009d7fdac;
mem[466] = 144'hf15009f8f9e2071bf6350061f964f184f013;
mem[467] = 144'h0908020407f0f6410de0080b03c0069a09bd;
mem[468] = 144'h0e5e00a0028ff181051e0586fe93ff06fb97;
mem[469] = 144'hf90f0f21fe1f0f6e0af5051a0f3bf6c40019;
mem[470] = 144'h0a89f0d5fe3c07c40aa7f31901c7fc6d0ba0;
mem[471] = 144'h0293f115006df590f317fa600e8c06c00b61;
mem[472] = 144'hfa420b560552f23ef59c03070a90faa2fe61;
mem[473] = 144'hf04503b0f420f7f8fc23f03bf117fbcafbac;
mem[474] = 144'hf0d4faca014304300dc5f477f3bb0b38f64d;
mem[475] = 144'h07b3f398fbc3052b05db09150022f598fecf;
mem[476] = 144'h0455f23ef379fd71efb405c70aeafdf5f598;
mem[477] = 144'hfb4c0f00fa2ff761ff67f23dfcbb0bfe0867;
mem[478] = 144'hfb0a00b50e9f0879f9a4047efa2ef631fbb9;
mem[479] = 144'h0a5ffecbf2660398f1520a8bf3200f2af869;
mem[480] = 144'h0c02049bf23e064406440f74f2dbfec7f452;
mem[481] = 144'h06290babf812086cfaef095e02240f850758;
mem[482] = 144'hf665fe330a6ff114f7adf0d00a3ffbb0f297;
mem[483] = 144'hfdde0ecaf42409b404d2011f0338fb540077;
mem[484] = 144'h04c60a59fab504760520f1540b8afe9c032a;
mem[485] = 144'h02290e34f874fb3af4f1ff85f3490925f5eb;
mem[486] = 144'h060bf4fe09ecf5f70d8e0250fdf9fc9500ab;
mem[487] = 144'hfe930fb7fad1f83df036f10ef10df2d409ea;
mem[488] = 144'hfa180e660f8104710f0bf7d8057aff3af43c;
mem[489] = 144'hf55b04c50822fdfa0313fbc2ff390e9bf878;
mem[490] = 144'hf6a206ed0bc1fd44f63f064ef38608befc5f;
mem[491] = 144'h0d6805ccf416f9a0f7de0d710a82f449f91d;
mem[492] = 144'hf400f6610f23f0b7f8f2088cfc3801060572;
mem[493] = 144'hfc1a012a07eff2a601a1037e0e05fa56f638;
mem[494] = 144'h0f28f3f70af60f1c0af40c76042a0a50f7b1;
mem[495] = 144'hfeeaf418f48afea20007fd5bf31e0423076b;
mem[496] = 144'h0a83f6de020b030bf6e6ffa4f810f8e5f961;
mem[497] = 144'h0e590412fdbb0b94f082f245f056016ef2db;
mem[498] = 144'hfe6ef1dcfd390b2e0223f73ff4610892f481;
mem[499] = 144'h013202f2f1c7fc43fe88ffb30c9cf23ff959;
mem[500] = 144'h05f9002104f60199f3f00c8ff9650483020c;
mem[501] = 144'h03ccfe3f0c57f6c20b4cf794f6dcf4940853;
mem[502] = 144'hf5480d4e092708bc0285fcb8fb270725f986;
mem[503] = 144'h0ce1f4b1f352f861f53bf48509eceefef21f;
mem[504] = 144'hfc54f28d02b7058bf905f6430215ff640dd6;
mem[505] = 144'h0403092304f5f2ea023e0c99ef1cf010f85d;
mem[506] = 144'hf0b50593fb3c038a0542fdcdf628f055f354;
mem[507] = 144'h07580a25f163febd0c500aeff867fd73fcde;
mem[508] = 144'h0a34f4690606fa98f3ec0632f5c9faf7f422;
mem[509] = 144'hf1bcfae20dba05360ae5fc9605a8f3ecf178;
mem[510] = 144'h00a303900b1809b8f375f55bfebdfd57031b;
mem[511] = 144'hfd57f42c09c4f156f76f0d36f5f7f7c2f14a;
mem[512] = 144'hfc0ef781007c0d52034800590d4af0f40cad;
mem[513] = 144'hfd2f0b46f209fde5ee790deff369f22c01ac;
mem[514] = 144'hfac003dcf2fb0dbf0377f8c5f7b8f222f8e0;
mem[515] = 144'h0d670d42fdee06c3fcbf045308cdfeb808dc;
mem[516] = 144'hf9b6fd61f6690e57ff200ab8f4640ac0ff56;
mem[517] = 144'hf4f3ff7108eefe40093ffb7100c1f07a0d5f;
mem[518] = 144'hfc63f2f30c3df58d036ef7d6f640097bfd87;
mem[519] = 144'hfce2f632fc3102f2061f02d2fda709b3f533;
mem[520] = 144'hf6830eec0a8df3070af0f18af9a40bebffc3;
mem[521] = 144'h09830148fdcaf474f7a90855f127fcd2f3fa;
mem[522] = 144'hfab50524faf2022df8aaf4830ad9fd7ef083;
mem[523] = 144'h05f1050c036af94a0005fdd7f932f1120377;
mem[524] = 144'h0a50f9baf01a0a450178fa140641f894f0a5;
mem[525] = 144'h0e7af9ee0205fe2401ddf517f4d8f76efba9;
mem[526] = 144'h0c3df8d502d2f9c00c4af75efbb0fc42f6a4;
mem[527] = 144'hfa320fa0f1e9039805f30f0304d20849f8a2;
mem[528] = 144'h0e8ef549ff640919ff140d9cfc0af3290e91;
mem[529] = 144'hfdd7fb54f103febaffb5043ef1900217f66b;
mem[530] = 144'hfcd9f8d9fb39036b03e90adcf790fefc0e27;
mem[531] = 144'hfc5df3e3010a0040f5b9018df17b020e00f9;
mem[532] = 144'h08b7f17c01a508a90b1803a5038ff743077b;
mem[533] = 144'hfb6402530e35fb140604fd31f490f7f6f9ae;
mem[534] = 144'h0269f1ca0ee60e4ff577081b0eedf2c2f4d1;
mem[535] = 144'hf906fda5f97b0c8d0f78004f02d5099fff2e;
mem[536] = 144'hfb520eb4f3a007abfb6c042df0ddfcc9f064;
mem[537] = 144'hfaef080ff8a6f74406c1096ffe94f46f01f3;
mem[538] = 144'h0a7f03ebf3010c5dff8100e505ca0e63f482;
mem[539] = 144'h0c6cfd94f5bf020df7a2f086f9c7fb920556;
mem[540] = 144'hfdfdfe8ff878fa2105e80978fdcbf79d0413;
mem[541] = 144'h05a6f6ce02970a40ff53f39c076a0ba0f2d8;
mem[542] = 144'h06e201500cc3057cff8b0cfe06d8069ffd46;
mem[543] = 144'hf0ae086af39a08d30d4df8030dd90c7a04b7;
mem[544] = 144'hf69ef472ff2b080d0944efc207d2fc4e041f;
mem[545] = 144'hfaf70a04f8930e81076c0adc0182040b0796;
mem[546] = 144'hfcd8fe10ff2bfed8f9020e5cfc4cf9cd0e4b;
mem[547] = 144'hfa18f5b8f06601e50e02084cfc220b9bfd88;
mem[548] = 144'h0795fca5f4550c8ff0be0b570b600cf3fa8a;
mem[549] = 144'h059bf20af801f6b30cc0f65902c30d06058c;
mem[550] = 144'hfbe30777f58f0a73f7b1f0940bf1f755fd88;
mem[551] = 144'hf173f6b4f3260a9e09adf72af0f5ffb80006;
mem[552] = 144'h0e0ef3a50d8efc0c093202b1f945f59fffc9;
mem[553] = 144'hf2bd0704f0c3f448fa6f0759098c06f3f54f;
mem[554] = 144'h03dff1f1f3210bef0b45f519f50ff1cc0d0a;
mem[555] = 144'h0e580ce2013b089906c901e40f61f635f3c1;
mem[556] = 144'hfcca06fefa20f25d0d10011405eefad2026d;
mem[557] = 144'hfc9e03a70b8bf99bf5c2f52200c6f2f908eb;
mem[558] = 144'hf2c803a500230a8af6e8fcfef6fe0af9f5b7;
mem[559] = 144'h07b103cbfb80087df9620267f0c5f69f0c78;
mem[560] = 144'h0827ff60f120080b091e0e7702e90b010b4f;
mem[561] = 144'hf7100cba09fc04ccfbe3fe9cf847f7f40143;
mem[562] = 144'h0a510e6e057ef08ff644f0dc07ac0897f0b2;
mem[563] = 144'h0437f65004d50700041bf0830b4b016eff3a;
mem[564] = 144'hfda40d74056407de002c060b0098fdcc00b0;
mem[565] = 144'hf08cfd670bd00c84ff900c29f4daf4f805d1;
mem[566] = 144'hff30f58a0983ff450f14073f0c050629f0e2;
mem[567] = 144'hf94a09cdf9710b2ef1e8008804d30b080ade;
mem[568] = 144'h0d97076f07bc0d4a04bf0afe0bf7f854048b;
mem[569] = 144'h0a550dc8fba6fb2bfba90be2f1bd0a4b076d;
mem[570] = 144'h0fd4f88709b1f30bf9ff01a80f1ef49bf8f8;
mem[571] = 144'h0dd7f9a0f6a0048b009effef09f70af9fc02;
mem[572] = 144'h02a6f17df442f591ffdbf127008101c0045f;
mem[573] = 144'hf6f804830e9a0697f907fbe00688f6e3fb54;
mem[574] = 144'h0750035ef09e08e3039d016ffbe40d240f87;
mem[575] = 144'hf88df1ab09e40b9bf8a9004ffc060d5cff2b;
mem[576] = 144'h0457fa32059efe340c39f290fd2c02870d9d;
mem[577] = 144'h01c2fe5effb5f85bf4670dac0a830ce90141;
mem[578] = 144'hf89bf28bfa64f9bf078508cffe26079709d0;
mem[579] = 144'h0e60f9b2fdd5fdf50647073cf02cfd72f8d4;
mem[580] = 144'h038e01230ced0cba082a041a09d6f75e0d58;
mem[581] = 144'h0ed6faeffbc10463038102b10217fe3af7b0;
mem[582] = 144'hf24f09c30c3ff5a3f4d90cb40760faf4ff98;
mem[583] = 144'hf5cd0eb40b6ff54b0458fef3f659f72cefd4;
mem[584] = 144'h0421fedcf84d0b53057603610bb0fd550573;
mem[585] = 144'hf920f300f10706d7f6dbefdf041bf50ffa49;
mem[586] = 144'h081afb8df2e5f764052df3c303e705a50ca0;
mem[587] = 144'hf5edf4140136fd030bba079efe5afb9f0de3;
mem[588] = 144'hfc0ff70406ef0b110edf05d6f31bf878f415;
mem[589] = 144'h0c540893f52bf482f1a7ffd9fbed03c507a6;
mem[590] = 144'h0760efdd0006ff160f02f9d104120dfd0ba3;
mem[591] = 144'h046f0964044008ea08dbfcfef4d7f34cfe9e;
mem[592] = 144'hf9870d4bfa4cf961fb23f42703290e09008f;
mem[593] = 144'h07b3f8aaf07c08c0fc93021c052dfafb03f5;
mem[594] = 144'hf61dfebe00d808c60e4efcaaf525fbc6061d;
mem[595] = 144'h0e2ef43800c00aeaeffa0019fa520ad7014d;
mem[596] = 144'h069dfd4ef1fb08fb07a6019efd74f60e0413;
mem[597] = 144'h07eef946f8430b9cf08d09f901ba0bf4064e;
mem[598] = 144'h0bde0e04f8b60b130d05043b04f30d27f100;
mem[599] = 144'h089ef7bd05790c93079f0b27fa25fa8df0b3;
mem[600] = 144'hf8b2007bffb6f0cf09fe01500de7ff6c063a;
mem[601] = 144'h00abffd3fad505da00f1f844f42af213fa06;
mem[602] = 144'hfa3ff776fae4f511f5f8fe840bb4f414fa3e;
mem[603] = 144'h01850ab20b1dfd2bfd41019c0df6f73efed0;
mem[604] = 144'h0792f7db0d1f0a230eac0002f140ff39fe11;
mem[605] = 144'h02fbf921038002a70bf8f0f2f1b0f548042a;
mem[606] = 144'h0644013905b1f9f605c9fda70290fc1a0710;
mem[607] = 144'hf7b7f619f65af4d50846f194f93b0ac1f791;
mem[608] = 144'h068506950d37f701fd640115f719fcd1f595;
mem[609] = 144'hf048f64a0ec4ef20f52f03f3fc51f588fe37;
mem[610] = 144'hf552fa34fd75fea30566f097077202c20f8c;
mem[611] = 144'hfd22078ffa5afd960888fc4b07f1f70203cc;
mem[612] = 144'hfed10287f2f3fcecf61bff20fb830dc30a48;
mem[613] = 144'hfd470632f3c8fcd5f961098e0d6208ccf355;
mem[614] = 144'h01f0f5be06e5fd67f779037dfaaf0b8bf43e;
mem[615] = 144'hfd4ff7540e2bf6160723f3d200d1f937fce9;
mem[616] = 144'h03e90af40b4d00830988fc050d58003d0c68;
mem[617] = 144'hfc5cffbc0f60faf9000602e4f2c708a6fd55;
mem[618] = 144'hf995f179f434f6a30bff0b8aefc302fc062d;
mem[619] = 144'hf82ef490053801010aa500640c550cd40be4;
mem[620] = 144'hfdeaf47ff3ce0ba70ece0228fa7c0d22fb3c;
mem[621] = 144'hfbc9f5070a260c00f814fd1fffad0d8106c7;
mem[622] = 144'hf4b90c5af755fbc5f3090554fd1504b2ef1d;
mem[623] = 144'hf59f0719f18b0b08f4d70ecff0ac04c902ba;
mem[624] = 144'hfc660656f15af8a10c81f605f572effb06dd;
mem[625] = 144'hf27b05def5fc0e68ff98f82cff5dfa03f08c;
mem[626] = 144'hf5ac0b9d014f093602eff400fab20531f2f7;
mem[627] = 144'hfb6cf25efbd60e12f490f7290182face0dd4;
mem[628] = 144'h0c790b5100b6fd31fa93fbab0467080a03ac;
mem[629] = 144'hf9e20b4204d4f1a10c3cf2ec04abf1870f9a;
mem[630] = 144'hf00b08b0f234f1dcf822fa1ef5360615f1d5;
mem[631] = 144'h090ef446f1e601200d8bfdcdfe1ef139f26c;
mem[632] = 144'h07df07910744f5cef70204360dd904cefe0f;
mem[633] = 144'h00a20c45f948f12df0e6f9bef68e00430884;
mem[634] = 144'hf5ba045d06860e04fc6cf250f5ab0b960f62;
mem[635] = 144'hf843fbb5f5bc0ecaf19b0528fb5c0283f44e;
mem[636] = 144'hff55073600aa06aa02fdf11001f8089bfb6c;
mem[637] = 144'h041dfd33ef440102fed7086ff5ccf78bf338;
mem[638] = 144'hf08d098dfe29ff18f4d4f5f101db0e16f09c;
mem[639] = 144'hf03ef16a0924f6a505ecf8d2f05a035efc2d;
mem[640] = 144'hf81ffce507720e550e4507b3f4d10460fcfd;
mem[641] = 144'hf06d0ac2053107b400b9043a072e05dcfe92;
mem[642] = 144'hf4f0f716fb47fac7043df035fdfdfe00f20e;
mem[643] = 144'h0f9cf5ea0018f3af08740f4af4dfffbf0d98;
mem[644] = 144'hf590feea0457045e05affc50fae50e2e014e;
mem[645] = 144'h019dff30f09af119f0030844f9f4f6e8f2a1;
mem[646] = 144'hf016fd130c2c04c400eef620eff6ffd6ffc6;
mem[647] = 144'h03d9010df40cf1dffacc0a3bf17df53ff54f;
mem[648] = 144'h0a78fc730ad2f2d60c23fb53f92df6f10261;
mem[649] = 144'h00a708eaf190024df8cbfbbcfc540dbc082d;
mem[650] = 144'h0dedf856f12ff0b80fc2fa3bf7b60f55f4eb;
mem[651] = 144'h0fc9fce407cef9e8f6f5f0650b690c450f42;
mem[652] = 144'h0b9002f1f25bf1b7fccefd91052bf1890aaf;
mem[653] = 144'hf54efb7802920c930bd60347f25f0df90583;
mem[654] = 144'h04fe0016014808590c3ff40b05920eab0dc3;
mem[655] = 144'hf96a046ffdf8f99cfd8df6250e96012dfa24;
mem[656] = 144'hf9eaf05a01f50f7806a9f7390468febffa97;
mem[657] = 144'h08fef00bf7030eca02d1f4990288f53ef6e8;
mem[658] = 144'h0f1607fdf6b0071cf7970798f420fe2b0a77;
mem[659] = 144'hf270f98208da00590373fa2df64efa960d02;
mem[660] = 144'hf50f0bf30d860996f489fa06f89efa66f330;
mem[661] = 144'h0ea70407f4c8fcee0564fc93fc9cf5e808fc;
mem[662] = 144'h0697fce90a28f57af7dff789f05203b90a38;
mem[663] = 144'h08c0079e02560c300cc4f5810d20fbc1f4cd;
mem[664] = 144'h094a0dc5fea3f7eefb2304aef0290809f0ba;
mem[665] = 144'hf2790a330a88f12c0066f2580b050fdefb49;
mem[666] = 144'h013df9a6f85f06430787fd5f027bfa1600c3;
mem[667] = 144'hfa7e05170d96f2f901a005490f190881f719;
mem[668] = 144'h0b27f1c5049e0d3d083ff34bf08bf004f466;
mem[669] = 144'hfc7707c402d0fbcdef030aa8f6e000fbf5cd;
mem[670] = 144'h05aef7cc0cc40dfb087ffe6efc9909f2f7d4;
mem[671] = 144'hf08af26bf6f906eef3ac0c06f0a80072f59c;
mem[672] = 144'h0aa8fea4f783f21f0b26f46c027af3b1f4b3;
mem[673] = 144'hfa730c88ff40f9ddfb54f00804e20a78f999;
mem[674] = 144'hf03f070df900fec3f429f68dfaaff101f9bc;
mem[675] = 144'hf89507a8fd8df3a2fab8f983f3d5fe40f7b3;
mem[676] = 144'hf18d08f406b506ed0096fc72f3ba08eeffea;
mem[677] = 144'h0b72f4f40b8b065cf54df31cfaee093f0246;
mem[678] = 144'h0285f83c0db30f7ef3c2f8a7f230fa4f09f4;
mem[679] = 144'hfad6f1bd06e904b707f900a2efbff211027d;
mem[680] = 144'hfb710825f0dcf0edf6dcf5b100d0f2ab03ad;
mem[681] = 144'hff180171f399f53f00f00f04036a0ad40119;
mem[682] = 144'hfe870d7502890469f28bfedef4f20441fdd9;
mem[683] = 144'h0a5a0cc6fafcfde30cf1fe27f218fe870a23;
mem[684] = 144'h000f05f70e6bf512fe7ff45f07ea04d5fb19;
mem[685] = 144'h08e20cddf28ff9270b84f00b0b600082fa6a;
mem[686] = 144'h0d3c02daf63ef3af0044ef5bfa71076f0260;
mem[687] = 144'h0f8cf0640667f7adf985ffbf04b50ca60f39;
mem[688] = 144'h0694035aff5d0d58047cf4fc0b2b0e6c099a;
mem[689] = 144'hfc5503710e57f8340a210988f6930f78fcfc;
mem[690] = 144'h0c0c09f701c6f66605f4097afef1f1780eb4;
mem[691] = 144'h07a5029dfe5afe600dc5f00df0260511fa60;
mem[692] = 144'hf97d01890cec0fe003a4f81a07a7f7ac0e0d;
mem[693] = 144'hf932f1b3fa29f3faf15a0fb302e400acf725;
mem[694] = 144'h03f301560993f969f6e9041307ac053df4c8;
mem[695] = 144'h024af8150cc8089803b70bcb00effea20a1a;
mem[696] = 144'h02cffbf30cd709ba0b17fde2017b0ed800e4;
mem[697] = 144'hfc500d380a9afb5ff9cc08a30984f41ffa35;
mem[698] = 144'h054208e90b630440ff130000f8530a8a0bed;
mem[699] = 144'h0da103eafe3efa5efbc90c8f0795042eff46;
mem[700] = 144'h09350b490b4800aa0a05fd64f307f31afa00;
mem[701] = 144'hfd8002660e47fe2afcf40dfaf304eff9fcc9;
mem[702] = 144'hf8c8fd6d07bcfec3f1acf1790229047902e5;
mem[703] = 144'h07e5082e0b0cf2c0f774f436fb660faa08fc;
mem[704] = 144'h0bcbff55f55ef5e70b71fbca04dff397fc2c;
mem[705] = 144'h0aa3f703f44a0fcef5320c630d250ead02e8;
mem[706] = 144'hf4abf5c204280c8f0f16f4390291028d0603;
mem[707] = 144'h0f8300bef88dfabe093a029bff90035505c9;
mem[708] = 144'hfa7f0324f5dff3c008d6f6baf9ce0487f4e2;
mem[709] = 144'h0be504f7fea901f5f9ea0552032af10907c7;
mem[710] = 144'h06de026ffd52037cfef3fd33ff47fe57052b;
mem[711] = 144'hf1430d9704fff665fa8c073ffb27f2ef06bc;
mem[712] = 144'hfdbef78601adfad507040888029bf4da03ba;
mem[713] = 144'h0d24fda1feda0fa908b3f4a90115f283fd24;
mem[714] = 144'h0eadf6b0f749044a01fd0dccf67703f9fff6;
mem[715] = 144'hfb460a59fe73000cf021fd1bf9d4f42d09b2;
mem[716] = 144'hf4c70371f452f03df7dff9bbfd1dfcaf07b2;
mem[717] = 144'h0cc5f5e9f02c0cb5f5ab003ef8a00a8c0bb9;
mem[718] = 144'h00c3f61809bb0c4ff1760c4e0c27efecf11b;
mem[719] = 144'hfb83f6e9ff8906850d2a09c30aa10e200f91;
mem[720] = 144'hf5380fb20286f784ffd0fa9801370724006e;
mem[721] = 144'h0130f740f22aff22fa44f6530f10fa54f5b9;
mem[722] = 144'hff14f34506d2f76d09510efff86401c1fa51;
mem[723] = 144'h0ed40c67f3670103f5d4f240f78df34e038d;
mem[724] = 144'h0c7b0c7efd0b0228f27cf0b2f78303d907c9;
mem[725] = 144'hf7fcfcaefa0ef506f526027b06f6f8e80b6d;
mem[726] = 144'h01450809f5a2f6a1fb6ffa5af8e4f84b0ab7;
mem[727] = 144'h0efff2c0f1320d43f66702ff0bc10c3ef7f3;
mem[728] = 144'hf1a50e3ef85dfa0b04fff911fda508defaf5;
mem[729] = 144'h0a76fa20face07ef023af63cf469f299ff91;
mem[730] = 144'h07ac0f54098cf7e003e00a71feb1fcabf5a9;
mem[731] = 144'h0b930697fbdf0664f9fff695080df9ff0b38;
mem[732] = 144'hf9aa0d330398ff620e74f1e3f4f9fbe808dc;
mem[733] = 144'h0bd4043bf14c0a52f986f22a0174ffff0067;
mem[734] = 144'h092109e208dcf4c1fe73f10ffe5604b5f6b9;
mem[735] = 144'hffe308a50cd3f7c8091409cc048a037e0a6b;
mem[736] = 144'h0bb4f252083101d3001f05d40d240f5e0c51;
mem[737] = 144'hf113faf1f252ff14f9e5fa0bf850f371fd16;
mem[738] = 144'h0d3b0ad8062304b904db00eb07e00b98fea2;
mem[739] = 144'hf338fc13f1fb06080c03f05d0abbfd1ef455;
mem[740] = 144'hf5f9f454f16a02b4fb9df0a5fc9d01c1fa90;
mem[741] = 144'h070c019a0884f6da03580e330704fae20551;
mem[742] = 144'hf562044d0a0ef9f8f5c9011cf1c4063cfd73;
mem[743] = 144'h0095060cf01c0b21fc15f728efdb0cfc049c;
mem[744] = 144'h0b4bfa94f503ffaf026f069904620101f045;
mem[745] = 144'hf2d5f57af80dfa13093d05e80c880d5b0791;
mem[746] = 144'h05a6f5b1f069f6a70d7cf601ffe8f090fc1d;
mem[747] = 144'h0544fe7ffc26fd8ef4070ae9f92cf6c309b0;
mem[748] = 144'hf448fb0201b8fb090b9e02f5fe14f7210a62;
mem[749] = 144'hf5acf081012d079902df0279f6b90375fb85;
mem[750] = 144'h018605fff2410423f638fe22feb8fe73f3d0;
mem[751] = 144'hf02cf50807fef86900b9f2320299febafad3;
mem[752] = 144'hfaabff5f077ef7510e050e85f83ef655ff39;
mem[753] = 144'hf189f244f9b3fe4af4bcf433ffa0f5d7f0ef;
mem[754] = 144'hff380bcef5eafd450766081e020400c9002d;
mem[755] = 144'hf791f974f350022404c8098904790313074a;
mem[756] = 144'hfdeff8c50feffa73003d0e2c038608700275;
mem[757] = 144'hf581f16eff54090d0e340e36032404d8f420;
mem[758] = 144'h0d4b03a20b1f05b0012e02bdf01cfdcef619;
mem[759] = 144'h06360417ffd3fac6f4f3001efd68f7840f2b;
mem[760] = 144'hff70feb108f50f21016503edfb880fcf02e3;
mem[761] = 144'hefa20c8405e60fbb03f8f51c0be6f7e40852;
mem[762] = 144'hfabef7b80f9108be087c00240e1efce3f9dc;
mem[763] = 144'hf18103d801a4f7e20528f891017bf786f3ac;
mem[764] = 144'h0b300e75099af12bf87b09bd03e60aabf048;
mem[765] = 144'h0c67fffef98507c606290819f9be0f3af86d;
mem[766] = 144'hf7fafc99ff8c09a40867efd80b3f0e790abe;
mem[767] = 144'h07b70f9807790783f485fc940b30f241fdda;
mem[768] = 144'h06f4feeeff2f08440e7af78c05b3f8d00703;
mem[769] = 144'h0886fa500aa603ca0acff8d1fa43f52d042f;
mem[770] = 144'hfe1ef4ef073b04edf5bffa330429f1f7003d;
mem[771] = 144'hfde0fb5b01d8feddf08df5d702820c34ef64;
mem[772] = 144'hfcebff68066d0fe4014cf8b3f39406960f4c;
mem[773] = 144'h040bf2b9faebf911f002ffb6f842f73c0cb4;
mem[774] = 144'hf611021c0aa2f35ffb68fdcbfaa5fc740cab;
mem[775] = 144'hf01807f203900f64efdbf7a6f9ef084004a0;
mem[776] = 144'hff5508ae066501bc0ca5f47ff5aa0a480667;
mem[777] = 144'h0a4304270fecfb58f1e204a4ffc80931fdf3;
mem[778] = 144'hf07c04890cbefdb8f5190c440d0a09d50b92;
mem[779] = 144'h00330e600ac20d97f297fe14fb9cfbda07b2;
mem[780] = 144'h01f5065503450083f3baf5aef31afe99fd23;
mem[781] = 144'hfcdc07b9f070f5c4fd34014ffc63f2b8efa7;
mem[782] = 144'h053afc04fc000a2ef1550331071e021cf870;
mem[783] = 144'hf257fa19f6520f1ff655f1b5fc080581f955;
mem[784] = 144'h09c8066d0b280c9c0347032af50ff64a0ae1;
mem[785] = 144'hf0b50273f357f9e305de0504005a0bf6092a;
mem[786] = 144'h0f9af05e0ee4fba10516054e0ba40b5405b2;
mem[787] = 144'h085ffef203ff0127fe60f9dafda502e202a0;
mem[788] = 144'h00cb02da0af8f7adf6d2062e05100846f40d;
mem[789] = 144'hfea7066202efff26fb37fa1101010ac90c70;
mem[790] = 144'h0c6bf849f55b02daf037fa72f025fa33f7d4;
mem[791] = 144'hf14000ab03b6ffb7fb7f04f4fdcdf7620d0a;
mem[792] = 144'h02a1f0740003060c029e03fef8e7fd4df477;
mem[793] = 144'hf5d8fb8c06ed079c05f10e05f64f077c0822;
mem[794] = 144'hf1bdf4ab05cefde6fbb6f12d0376f9230c56;
mem[795] = 144'hf2520596f47cf2320967f87a00cdfad202d9;
mem[796] = 144'h0ac104ebfcb204b805a9072f069d04cf0ce8;
mem[797] = 144'hf319f11901cbff8cf7950432f10ef7dc03f1;
mem[798] = 144'hf9bbf483fc39f2040a07ffde04cc0f5a0203;
mem[799] = 144'hfbea0e90f0b50a21fd8107570776061302fb;
mem[800] = 144'h02e3fd5efbb505abf0f2fa30f738020906de;
mem[801] = 144'h087f049ef64ef4a5018508490a6bfbb50e20;
mem[802] = 144'hf684f485f33bf44d04d2091305e106f3f0b1;
mem[803] = 144'hf69c060b05c2f62ef438fc64f00dfa67f398;
mem[804] = 144'h03350aee0e2702de0cfff904f54bff07f1d7;
mem[805] = 144'h010afb760ae8f0cff81b04c405c0f6b5001a;
mem[806] = 144'h0f7b034505b5060e08f2f0a408c4fb46f648;
mem[807] = 144'hf704ff85f6cef5ca090f03e80283f401fe58;
mem[808] = 144'h0c2bf9240ec0fb1ef9900139ef75f42e00a8;
mem[809] = 144'hf2adf5cbf3d8f8e609660e5f0bb6f64ff803;
mem[810] = 144'h05faf8dc069306df0732fb04f2acf02ef183;
mem[811] = 144'h074bf31df9590932079a0bc9f9bf0a58fb1d;
mem[812] = 144'hfc91f3b6f53d09ddf0140b640a430db7fb42;
mem[813] = 144'h04140ad507f90c0f0ee9f013fc51f44ff3e4;
mem[814] = 144'h0632ffaaf4480e55f6f1086e0cea0cc90f05;
mem[815] = 144'hf50df6980e650ba0f9200f17f99904b00027;
mem[816] = 144'hf8110855f8edf4f30a480d61f0a10a51fb3b;
mem[817] = 144'hfd670a270e84ef7209570682f93000ca07e2;
mem[818] = 144'hf0acfd560498f86205340d4bf2cb0342f0e6;
mem[819] = 144'h09adf903f8600c3af56df029f9bc05daf369;
mem[820] = 144'hffc300e00ae1f5c9f26a0c230c240a62f47b;
mem[821] = 144'hefebf855f1b4f193016b0dc40d5f026a069c;
mem[822] = 144'h03f2f89b06faff80ff12f8bc07c309dbf307;
mem[823] = 144'h0ac90ebb035b07860115f66ef072f5fef5f2;
mem[824] = 144'h01d70ca8f7ad0540f55d0b19f182fa990140;
mem[825] = 144'hf00df315f2a3f037fdd5fed5fc41f2e8fd14;
mem[826] = 144'h060208c600340c8ef861084806a60a24efb8;
mem[827] = 144'h0eea0781f9bef16bf6820dcff0bcfd4dff03;
mem[828] = 144'hf40f0e400e3cf3770212ef95efc608b504d8;
mem[829] = 144'h094cf89a0a570958f235f3af064506d7f1dc;
mem[830] = 144'hfa6dfe06fa1304cdfa28fbc3f7bbf5480116;
mem[831] = 144'hf0f40eecfc9400350fbaff130f0803e20ba3;
mem[832] = 144'hf84b014502f5f3e0f8e10ed70d2af16d0908;
mem[833] = 144'h0352f9ee0e25f5da02d5096407d7f16ef3f3;
mem[834] = 144'h01c70815f423f4f50a58028903fdff20f5e4;
mem[835] = 144'hf87c09de0755fdffff63f66c0addffb3f7cf;
mem[836] = 144'h008602b7f4dff0d9007e08670654020e0f93;
mem[837] = 144'hf757f27402bd05b0fbeb047f0685fbd1fb71;
mem[838] = 144'hf876f6bd081707c1f335fdd80394f7d1effd;
mem[839] = 144'hfb930dc405a30f8df75d003e0a3f03c8fb01;
mem[840] = 144'h030df04c0277f9b8027d0db7f8b6f271f379;
mem[841] = 144'h097efdb5f669f67d054afcaff77df51b0c0e;
mem[842] = 144'hf5bc022208bcfd12f2c002f0f7570e8bf080;
mem[843] = 144'h0b72f6a8f128f89efeaef105fea30375f28c;
mem[844] = 144'hfc2b03e6fa28f35d033af808ff0ef56b05ca;
mem[845] = 144'hfb80f490f70e0284f7d2f08efd68057f0009;
mem[846] = 144'hf030fcb40f4e092e0c7804fdfa16053ef753;
mem[847] = 144'h06650d900ef70f4107a9f7a9012afb880a1f;
mem[848] = 144'h0693f084f3c8f2e103eaf38ff26bf8faf3b7;
mem[849] = 144'hfedbf199029dfb13fb1c0434043a0842017d;
mem[850] = 144'h0238f29a06c802d60f64068a0f54faaaf921;
mem[851] = 144'h09f2fe870ebafab40086f925f2a3fbac013b;
mem[852] = 144'h09c00f3b07f5f7c4017ff088053bf2dbf573;
mem[853] = 144'hf923f1a20a32fa83f53aff6608ef09100571;
mem[854] = 144'hff97efac034404aafc680946f4d50332062e;
mem[855] = 144'hfb42f225fc2b03af0ea30a97f6e8f28f0f94;
mem[856] = 144'h05e6f20a038dfe7b0878fa47fe7ef3cdf6dd;
mem[857] = 144'hf5b8fc4ef8e1f8cd0dc702a107f5fa6108b2;
mem[858] = 144'hfdfffa600e35011df36b06c1ff690c6afd6a;
mem[859] = 144'h084aff7ff88705890bc4027c053e0ed4fcc7;
mem[860] = 144'hf6160a5602350e08f7d6f5150b1f0ce00642;
mem[861] = 144'h08e1f79307b9046509f307a809c7f213f003;
mem[862] = 144'h0e81fa54fff809600c73f7bf0ba4f496098c;
mem[863] = 144'h01c2fed30a1e00f30be7ffb801910fcb04b5;
mem[864] = 144'hf0c2f4fd09b604d2f4850183f650fa390e98;
mem[865] = 144'h00ccf36cf75dfa34f427f35b0e17fffdf8fb;
mem[866] = 144'h0ed802af0548eef0f86afcbcf28f03e5fc24;
mem[867] = 144'hf36100bf02ec0362ff000fadf8f4f6fdf13a;
mem[868] = 144'h09f8f24ff0bdf117f4d1fc760f3ff025fa3f;
mem[869] = 144'h02b3fd83f1c0f03700990139f2eef8f8ff2f;
mem[870] = 144'hf07afeb106470691fd12fcb7f6c1fc180b5d;
mem[871] = 144'h054bf4e1070109ec05b30d0304ca01630c01;
mem[872] = 144'h0d52f28bf1f5022508bdf1fcf51cfcf2efe8;
mem[873] = 144'hf30e09b30607f6c8094ef59a0a21f5b1fa4e;
mem[874] = 144'h07190052f8f0f337fb5800c6f2dff843f898;
mem[875] = 144'h04b6f6a80959f61605ab0d76f89b096d0bb9;
mem[876] = 144'hf75e0a71fc430f02f8c70490f839fea90cf4;
mem[877] = 144'h0f01f78c0a81f83ff4bc0c960bed0f31f966;
mem[878] = 144'hfa4a09fdfd830906ff540d990f1609e0f3b5;
mem[879] = 144'hfa860e1005ac0d950608f4a80722019f0228;
mem[880] = 144'h0e120539f2b3fcf405b708c6f7e10ece0959;
mem[881] = 144'h0272f0cb0034f0480d9afe06f307f51d027a;
mem[882] = 144'hfbd006390e830a250a87019cf2b1ffc4054b;
mem[883] = 144'h09a2f4d9042b0a1e00840a2f01440c63fb86;
mem[884] = 144'hf861f45f084bf87306a2f36dfede0f04f1f7;
mem[885] = 144'h069ff1950bd40ebc0a6df66906ebfff3f0d8;
mem[886] = 144'h0ee3f422fc910ce9f25805e7f9d9fda40583;
mem[887] = 144'hf9ea0702039e02c909e5f1dafab005860c38;
mem[888] = 144'hf4c8f44405580c2df0450947f943fb640ded;
mem[889] = 144'hff76f596fd6a095b0eb7052101780dc70a06;
mem[890] = 144'hf8a309f0f0230c1af3e2f4290858f2050d45;
mem[891] = 144'hf322074c0d90f07dff420f71f6def3d60f99;
mem[892] = 144'hffabf544f70806b4f45efda7051304fffddd;
mem[893] = 144'hf55f073d0ad2fc6fef72fbd00bc0f623f8a6;
mem[894] = 144'hf5e1016eef9ef26bf6baf26e025df7510c2a;
mem[895] = 144'h09f705b5067afcc7feff059a0ee7f927f424;
mem[896] = 144'hf09104f10e7901e300cafc04099106650015;
mem[897] = 144'h0eca0b79f023fc180b78f5ad0185fb0cf180;
mem[898] = 144'hfad6f1d7073c0686fc6d0e8c0744007a0b06;
mem[899] = 144'hf2eb085ff6b3fc54f0fbff790b6407bbf827;
mem[900] = 144'hffad02f1f51c0b49fce304fcf57df0af035e;
mem[901] = 144'h01ef0327f5c9026ffb530b40ff08fa5af3ea;
mem[902] = 144'h0d390f40f0ab0cfeff63fceef8de0feeff1b;
mem[903] = 144'hf7ecf76906570cbf0ca3f5370bb002cc043c;
mem[904] = 144'hf204fcad08a7033b087ff49ef0bcf646f3a6;
mem[905] = 144'h05cdfe6ef6f0fc7ef4870977013306ff086c;
mem[906] = 144'h0e3d0438fe4b0123f0c8fc64ffb60a79f4d0;
mem[907] = 144'hf2dffb0504ae05d4049cfeefffb4f0c4fd92;
mem[908] = 144'hf9900d23f32e03d307fc0b47f5d2efc8f529;
mem[909] = 144'hfaedf7260745f8c8f833fde9056ff5c20bc5;
mem[910] = 144'hf2aff309fbc70f35f78f040e0940030e0a84;
mem[911] = 144'h06bd0c400ac4f915fb48f41b0dfa00f5f131;
mem[912] = 144'hf1fbf3fffaf205f1086ffce9f0a60c8bfa17;
mem[913] = 144'h008ff12af0cd0f75f2a10efb0c64f65d097f;
mem[914] = 144'h0c15f5e3f21d03a1f388f0530a390ccb0ba2;
mem[915] = 144'h0707fe3907f0f9cef0170fcdf9260b6bfd19;
mem[916] = 144'h054003140af50db5f591005e03470f470276;
mem[917] = 144'hf02302a9f5c10db302360bf700f0f67ff90c;
mem[918] = 144'h0a92ff7a02ecff28efb4098b0b5ffe9f0957;
mem[919] = 144'h01acf8e0fe9bfa0d023c0ed50011f281035f;
mem[920] = 144'h062cfb35f4f9feb808be0f450b23f9a206f3;
mem[921] = 144'hf5e40279ff02fe050288ffd2fdcff5b30288;
mem[922] = 144'h051af929f649fb690948ef55feda0ec7f3a3;
mem[923] = 144'hf0b801fbf223f01bf53afb90ff9e05310623;
mem[924] = 144'hf796f3d804690d6c024407b6facc0e870544;
mem[925] = 144'hf2eaff67012202da0727f0f60af7f9e7f830;
mem[926] = 144'hf825f2d00f8d085a065efcbff585f50cf2fb;
mem[927] = 144'h037ef0f60a11070af2da0c03f88a053107a1;
mem[928] = 144'h016c095ff690fa990577003bf213016d0bcf;
mem[929] = 144'hfae9f1ed07610a720b24f7cd0067f31ffdd1;
mem[930] = 144'h02fcf5b2ff16fc9a039cfe99f43bfb23fe6f;
mem[931] = 144'hf933f744f1c50c370f13f4d20def04ce060c;
mem[932] = 144'hfce6094304160f45f5880968096a0018fadf;
mem[933] = 144'h018bfa9bf840077c019f0b5dfc08f50cf159;
mem[934] = 144'hf610f7ce042dfad1fb7e01450342fad902bd;
mem[935] = 144'hfc3a08f1f03708380341f061f49b0d84f9b4;
mem[936] = 144'h053ff94c06be047cf71cfba7f6ed0556f1df;
mem[937] = 144'h05a80186f4f404ac019404fef020f381fd65;
mem[938] = 144'h0fc2f1f6fdbbfded05eff965f19705c5fa16;
mem[939] = 144'hfde5f5d102ab0555f39af739f87007f0f154;
mem[940] = 144'h0ad9feeb0e5c018b09a2fcf1f7f5ef960170;
mem[941] = 144'hf730ffb30a18f18b059bf230088afae8fc85;
mem[942] = 144'h0b9cfb4d08caefe8f9d406a4085c0bf40ca9;
mem[943] = 144'hf54d0a0800070343f47b06faf71cfeb40e4c;
mem[944] = 144'h0ea80a500c4403e203380a550d0b0408f212;
mem[945] = 144'hf73af8c1fc35f37e02cf0ddb033defa0fb40;
mem[946] = 144'hf128fe9403eef4c50c970601033202e8f382;
mem[947] = 144'h0acdf05a093ff054f3f5fa96f4bc01d0f20d;
mem[948] = 144'hfff4f010fa3a0556ef650733f38d0cfcfddf;
mem[949] = 144'h0c03f94df4ce0ac5f8fd0cc0fa31f033f592;
mem[950] = 144'h04f80262f66ef6100974fca2faac099401fe;
mem[951] = 144'hf9c6fdb705c9068600a7f25103630a0e060c;
mem[952] = 144'h0516f809fbbef13a0b3e095cfe74ff0f0b54;
mem[953] = 144'h0c6d00660631f63e02c0f2e00ca003880441;
mem[954] = 144'hfd35f8d8f132002cf60bf89af17a0ba90752;
mem[955] = 144'hf7acffff019308a2063bf1dd05bd097a0db1;
mem[956] = 144'hfdf8f5cf063ffd670cd6fd70ff72f098032c;
mem[957] = 144'h0e01fef8006ff8e104b209410962fc9002d5;
mem[958] = 144'h0ae4f0b70e90fe7b0752f00c08ca087b03df;
mem[959] = 144'h0d150209f1900936fb96fd2e0934fddafd9a;
mem[960] = 144'hfa77f55004020c100496f3fa0ea1ff340afe;
mem[961] = 144'hfffbf1d8f1d309f5ee93fe87fe7ef977f1c6;
mem[962] = 144'hf8fcf5d6fdc50d8ffc73007005f3f6d2f701;
mem[963] = 144'hfc5c0d6f0967fef6fa8b0e69ff450144f62b;
mem[964] = 144'h05570e2d08ed0228f9b1fd36f292f85ff06e;
mem[965] = 144'hf426feaffc3f04b0f80d096e0113f68c06d2;
mem[966] = 144'hfa59f9f90dda090d0e94f20204b201d5028c;
mem[967] = 144'h0206075505410389fbaa0357f036f2d80090;
mem[968] = 144'h02e7f7b7f4e307360d200225f42cfe2c0d76;
mem[969] = 144'hf8adfe30fa2603bc04ac02e2f13d0a10f8a7;
mem[970] = 144'h0974f523fe3cfbdc07920b01f9000898fb7e;
mem[971] = 144'hf29afb5e0c84f3f8f9ff047afddafd7ff185;
mem[972] = 144'hef74072c0b1c0654f832f1fa0d87ff44f770;
mem[973] = 144'h070d05acf0cafcef0d080f89f1ae0a65000c;
mem[974] = 144'h0d8307bb0a98fa2af2f00acd024b011fff42;
mem[975] = 144'hf253f02fffc70ca3f79707af0c43f82ff77f;
mem[976] = 144'hff61099df7660e4ffb380ccc0d41f1c308c6;
mem[977] = 144'hf9e4fba9fc1c00a80e0e0c0e00c6fafa06a7;
mem[978] = 144'hfbd20c450aeff0b006cd057ef698041bf8ad;
mem[979] = 144'hf626f614f56ff8410a150f46014502f00a9a;
mem[980] = 144'h017401aef05ffb8604e10649f116f4b50903;
mem[981] = 144'h06c0089bf5cf0b930093027800dff0aa0ccb;
mem[982] = 144'h09830381fd380044f9c60b2ff4d0f358f036;
mem[983] = 144'h0e03f5de010c0c6c09dc0f8902d30d73f163;
mem[984] = 144'h036ffac403b00374f5b7fdd5f48901e3f832;
mem[985] = 144'hf1a500c1f6d6f83af6a409c703e007260a96;
mem[986] = 144'hfc0708210f56f71efa2df44a05c70607019e;
mem[987] = 144'h0ec1fc690baef741063c0fd10dec098e0447;
mem[988] = 144'h0cb70195f66d079e07c1f0c6fca5f9fa0f33;
mem[989] = 144'hf80ff74b0300f830f136f9d6fb58014ef2a7;
mem[990] = 144'hfec1f1eef4f80342fe9d01b30e26f30f0768;
mem[991] = 144'hf57efa3af458faf60d01fe3a0091fa790bd1;
mem[992] = 144'hf7250aeef3bc08300fe4f915f2c9035bf4e9;
mem[993] = 144'hfb08f05ff38c05f3fb460ebdf29c00200f84;
mem[994] = 144'hfc3bfe09fa09fc58f726fe0a0d01061dfbad;
mem[995] = 144'h0bfefdbd0ad4f440075ff849f77ff7a509c2;
mem[996] = 144'h0017f4b1fb5cf4e1f886010cfec2007a01d7;
mem[997] = 144'h09e9f7c8f629f6fe0c790152f09c025d0201;
mem[998] = 144'hffe6085a0850024ffe8f0b500c7c0a90fee6;
mem[999] = 144'h00810bf10cbefcd1f1200148091cf2440f2e;
mem[1000] = 144'h0375f6fcfd940c4e0f4afe39097af1310ba0;
mem[1001] = 144'h0bde060a0f5203b407d505910048f246f91a;
mem[1002] = 144'h063d00f4f4770abc0c92f606011d07a3f2e7;
mem[1003] = 144'hf592f51d03b3fe69faf0f721f3cbfe12fc99;
mem[1004] = 144'hf0af0b80fc520bc40ede07d30066fcbff4f5;
mem[1005] = 144'h015808120baff273f2d0fabc05c1001c0c82;
mem[1006] = 144'hfde70127012700e9f868f0befc5d0657f328;
mem[1007] = 144'hf0970a58fdd70aaaf1c6f0660b1ffba0f4d5;
mem[1008] = 144'hfd75f02505b80050f27bf2f6fd81f771fe70;
mem[1009] = 144'h07c1ff25f555f7f9fdfe0b5b0267f990075b;
mem[1010] = 144'hf4b1ff72fa000548f75ff6360d7c0cf8fa67;
mem[1011] = 144'h0db7fb34f99ff868f36e0d2cfcc8efd7f5a4;
mem[1012] = 144'h04f2fbc40594ff510be8f7a708320c6e0aa4;
mem[1013] = 144'h09c0f2c0ef22f941fab0f793f120f830f6a0;
mem[1014] = 144'h09c5f5730559f005f7ae090e0a40f2dceed2;
mem[1015] = 144'hf2310d100bfef1510ba60867f960fc6d0ef3;
mem[1016] = 144'hf14b099ff1ea01e90025f5450e1c0640077e;
mem[1017] = 144'hf6d1fb61fa41f497efe0f439fc4cff8506a0;
mem[1018] = 144'hf4ff03a9f379ffb001290594f88b006e06e5;
mem[1019] = 144'hf1a1f3620c5d0478faa5f7ea064c0051fe50;
mem[1020] = 144'hf802f6ba0c40f52ef2950d34000f0cd70a52;
mem[1021] = 144'hfa6902e70ae9042404f1f81af137fd18031a;
mem[1022] = 144'h00c6023e089ff374f56507e600dd04bafe0d;
mem[1023] = 144'h032e00040ecdfdc7059303050f91fefaf157;
mem[1024] = 144'h09a70a1105ce046ef220fbfdf9a60376f909;
mem[1025] = 144'hf19dfc410a6303ecfcd3fd06fca7f295efdc;
mem[1026] = 144'hf95df8b4fc2b0ed7fca9f116f902f9c0fbf1;
mem[1027] = 144'hf3cf04b6ff33f8ebfd4ff0c70006fa2bef89;
mem[1028] = 144'h0528024efd6af002010209a0f864f701072f;
mem[1029] = 144'h0796f94a09350aa7f636f727ffee05be0475;
mem[1030] = 144'h04cbf27aeef8f2bdfbeffabffcac0525f469;
mem[1031] = 144'h0e8601ce0309fcb70b79f7f4f2d8fc17ffbe;
mem[1032] = 144'hf3c307edf08ef7a3f5def685fc58f7bcfdd5;
mem[1033] = 144'h0776f158fe72ff6bf696fbac0681f419f1ed;
mem[1034] = 144'h0c700316fad708eefd4902d2f3e7f0d504ae;
mem[1035] = 144'h020d01c90b71f40408790d80098500940e6f;
mem[1036] = 144'h0b8605070a13036f03aff80ef169f9a3fa09;
mem[1037] = 144'hf54af098007bf9e20e0604d9fb81f23efee4;
mem[1038] = 144'h0d6f0ac7f44df7bbfa8f0356fe0500dbfb17;
mem[1039] = 144'h01e5fcf0fa0808b6feea038cf85e0495fa1b;
mem[1040] = 144'hfe45fa91fcf10597041c01a80953fdc1fb34;
mem[1041] = 144'h0de20d4df46b0cba0be8f07c0369fd43098e;
mem[1042] = 144'h0d5a020e0b40f3130c3cf7b3f439feb304c5;
mem[1043] = 144'h09f6fdacfca9f344f8aefede002aff080c2f;
mem[1044] = 144'h03750452f16c079bf9b206bd0595fcb2f990;
mem[1045] = 144'hf699fb3d0f26f7330384fd5cf6d904340cd7;
mem[1046] = 144'h04a30b0bfe4c06e2efe402e80a980a62fe30;
mem[1047] = 144'hfecbf3b0eff5fc3cfd900f4f0caefeb108a2;
mem[1048] = 144'h0f090185002ffef0093cf3ea0a7703d2f402;
mem[1049] = 144'hf3b9f9f8fb47f2abf33e05400045f5ecf86c;
mem[1050] = 144'h0824f5260d5eff4a09c8f9ed004e079d02cb;
mem[1051] = 144'hfacbf4070a3c022effb5f0700c0b0336fbb1;
mem[1052] = 144'hf644f491fed80731fe360af8f72b0b6c03ee;
mem[1053] = 144'h0eecf224f347fa7ef5c0f943fae6f03cf951;
mem[1054] = 144'hfdbdfc71f08ff18d0d47ffeffaf805a6fcc6;
mem[1055] = 144'h09f5f6110d87fb36f85ff9680f0e03dd0bc3;
mem[1056] = 144'h0d37fde70796f737fe11f4f8f42b0d2106d3;
mem[1057] = 144'h0d7bf248f136f088f02bf5370e970b2a0f89;
mem[1058] = 144'h0a7a0a36fd5a0df7015e08a1f626f54004ba;
mem[1059] = 144'hf48bfb1c078cf008fd9001cc00c009150edf;
mem[1060] = 144'hf7c1014afc4c02490519f184f6a0f13bfce2;
mem[1061] = 144'hf93b00f2fe0cf675f745f61dfc280d7ff635;
mem[1062] = 144'hfdc208cbf7b5f5b30653fd8afe51fa830346;
mem[1063] = 144'hfd0705d70b250f58f92c0011f233fad5f418;
mem[1064] = 144'hf4690d9dfe650d76f1c80da3fe84fafdf248;
mem[1065] = 144'hfdb4ff2cfbdb00cffaf1f6dd059702b7fb27;
mem[1066] = 144'hf2e3f25af8ebfd6ffd1af5750c0bf5d6f911;
mem[1067] = 144'hfa78f25f0cc0f3870d4405bf069af2a20e56;
mem[1068] = 144'hfc0ff90f09e4f4a7f2ccfc74f9fa078ef0e4;
mem[1069] = 144'h02a303110a8ef40dff06fb2a0a6afd5803c2;
mem[1070] = 144'hef83f647f9310d310094f388ffb90670ffa5;
mem[1071] = 144'h00d10309fb89f97bf08c0586fe52f3f60fa8;
mem[1072] = 144'hfb57fb3e03d6f5b5f786f9a4f2b8f7be01f5;
mem[1073] = 144'h0aca03560574f35c00fb0166f897036d0e33;
mem[1074] = 144'hf91df0e9fac3f624ff1defc5f25ef2380f96;
mem[1075] = 144'hff6708fef3af0f01fa31f0a20149f2f90a63;
mem[1076] = 144'h076dffa8f9b10783f656f0c1f0cc0200fec8;
mem[1077] = 144'h05940cd2f6bbf9cf0d9e0290f207f48cfd94;
mem[1078] = 144'h06670c770019f6ebf654f963f2e80f30055e;
mem[1079] = 144'hf6e90e33f047038102e6f7bb0d71f887f572;
mem[1080] = 144'hff5a098108aff4ab0c9400850593f2eff26a;
mem[1081] = 144'hfe3905def12300ccf17afadb08800e66f115;
mem[1082] = 144'hf84ff9400762082afe86fe2ef8fff8cf0231;
mem[1083] = 144'h08b00b460bc00f7d036f053ff8e60c190496;
mem[1084] = 144'hf73805a0ff79f50d04a00ab8f113f9cdf43b;
mem[1085] = 144'h0c8af0a002fdff9df7390973037c0b22053c;
mem[1086] = 144'hf989fcb107d8f8c401de0c860623079303f6;
mem[1087] = 144'h05800bfaf38709be04cafe0eff2aff0807d2;
mem[1088] = 144'h0c1205cd06d8054e01ccfbb70b2ffe9e004b;
mem[1089] = 144'hf9270982fe28f6fcf6710f0bf78400c9ffd8;
mem[1090] = 144'hf09afb23efb70d3a021ffde0029ff404f644;
mem[1091] = 144'h036bf7ea0c89fffefd77f8aff9bcf5080493;
mem[1092] = 144'h04d7f608fe3cfc1afe3cf35f02d9f17f03bb;
mem[1093] = 144'h028bf7e3044b0ac206940ed4fd9ff7690da8;
mem[1094] = 144'hf398efd50e38f60ff5cb001b02240c75fa45;
mem[1095] = 144'hf9bd083d0d17fda407ebfdff04e3f555003d;
mem[1096] = 144'h0bac0b7dfc6d03e60875f29af861ffa6f07c;
mem[1097] = 144'hfe50fffff3fef9c00adf04530a39f9b7f53c;
mem[1098] = 144'hf48700cff651f174056e052c00b00ec40b58;
mem[1099] = 144'hf1ec0481fcc904f411c6f64d0b99f8edf201;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule