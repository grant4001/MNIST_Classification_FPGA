`timescale 1ns/1ns

module wt_mem6 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'hffd1f06c10710259f4ebfd9bf12cf5a8097e;
mem[1] = 144'h0312002c0078f27506a8f75a0bea07e9092f;
mem[2] = 144'hfba1f652f8e40015077605760b630aaff868;
mem[3] = 144'hf1a708e70bdd0c6d035a0d210237fcd7f6c0;
mem[4] = 144'hef48ffd4051500fd05d007a800d5f005f96b;
mem[5] = 144'h080af471066d00daf0acf618faa1fa6b06ca;
mem[6] = 144'hfeff0c6ff6450af7052c0853f3500d0cf0cb;
mem[7] = 144'h00b1fac30733fbabfeadf28cf0aff6870d37;
mem[8] = 144'h07d606540692077c04f4f54cf57cf8250dbc;
mem[9] = 144'h04a3ef7cfb21fbbb0f42069f07eff0e2f74d;
mem[10] = 144'h071d0c4006e70a000f6c054f03d60855fcdf;
mem[11] = 144'hf59e05b70482f0aa0d5b000e00d9fc7d00c3;
mem[12] = 144'hf23ff8fe059af298fc76f932f233f2e7f8af;
mem[13] = 144'h05880123fc6107adfc7409ab0748f830fd74;
mem[14] = 144'h0539f4fd0997f31f0856f3fcf0870bca0ab7;
mem[15] = 144'h07d20675f71a0d1af461fcdffcda0749fb10;
mem[16] = 144'hef18f353fc4df94b0d8dfde6f2e90de0efc7;
mem[17] = 144'h0aaaf7aaf0d30c09ef1a015901790e46f445;
mem[18] = 144'h0af0ff63f981056103d80c17f1f80eb00546;
mem[19] = 144'h08f2fe600d3cfd2cf9b90bd30649fd26fd2b;
mem[20] = 144'h0cfc0dc9022c06d7fc8fefbb034af8e5fbd1;
mem[21] = 144'hf16c0b950ba0f8b709f1fc5df80b040bf8e8;
mem[22] = 144'h0d57f96ffbf0f52005a30713fc8d0d810a44;
mem[23] = 144'hfa06f7a8046e00820a300371fa22fd7dfc3a;
mem[24] = 144'h05fffea5eeca0c07028df8d0f19e03aefe50;
mem[25] = 144'hfb1f030c0cb5f030fb820a43ee92018aff87;
mem[26] = 144'hf11efb2b00dbf819064408befbdc02edfb0e;
mem[27] = 144'h0352f91d03a206590755efbdf35a09aef053;
mem[28] = 144'hfde40b46f7520ad3fcfd02050d3ef48afff6;
mem[29] = 144'hf254f3ddf91bfe3cff95032606a200740f2c;
mem[30] = 144'h09daf871f60e0040030c0de9075ef57c0335;
mem[31] = 144'h028ff1d6fa0a0d0a0791fd21f04202e0fa77;
mem[32] = 144'h0ac008ab08bf085f026b0998fbc60d05ff07;
mem[33] = 144'h07c9051308490f22052f0cf5000aeee0ffcd;
mem[34] = 144'hfcdcf1c203c9006b04c6ff6806c8044cf062;
mem[35] = 144'hf344f54605a6001b039d04cbfeb7fc02050b;
mem[36] = 144'h04630210087604df0761f5dafe9ef33f0f48;
mem[37] = 144'hf5d507c6fae5fc57fc470f81f3e9017dfc59;
mem[38] = 144'h06d4fd31f2e2fabbf8b60066f3b7ef3ffce8;
mem[39] = 144'h0995044dfcd20f08f64ef8080377067cf583;
mem[40] = 144'hfcdaff42f2f20e3cf72e0db2feca0051fffc;
mem[41] = 144'hfceafe48080b087effd6f6e7ffe2ee5100be;
mem[42] = 144'hf6dc039a08300147f429f4d2efa50ae2f470;
mem[43] = 144'h0b050bf106040cd0f735fc84085df3000433;
mem[44] = 144'hfce4f142fcba0a2bfc220ebff822fbbe0eb0;
mem[45] = 144'h02edf0cc079f02a80836fe9a0b090d43fb3e;
mem[46] = 144'h09d4ff0df9920e0e094df1f6f9b8eff40a1e;
mem[47] = 144'hfd7c08ad0249f88e01d2092bfdcd08a01077;
mem[48] = 144'h0ccaf9aaf960f7450dd50b0af9e40316f33d;
mem[49] = 144'hffc5f7170a3e00c1ffbd07f00a82ff730411;
mem[50] = 144'hf1ff008409780a44f1b3f756fc09f34d0d11;
mem[51] = 144'h047209e6fc2b064c015afba5fc80f542fc4a;
mem[52] = 144'h0e0304dffe21f83f054cfb9a0c040a91f1a5;
mem[53] = 144'hff88f4fa064df7f8074b0bf7fe7cff2302d2;
mem[54] = 144'hf162fa52fb190d88ff8bf658f6a4056f0a45;
mem[55] = 144'hf4bff9930648f1e4f2f3f5e70e4bf5a1f76c;
mem[56] = 144'h0750f6e306c6feddf467fac0f708fd85f3a5;
mem[57] = 144'h0bb30d1e0abb0e38f530f0a9fdd1f08e093b;
mem[58] = 144'hf1f00b57fe1e040bf7cb096d0ba201760062;
mem[59] = 144'hee8e091cf78ef0f7ff83f914ff35faf7f50a;
mem[60] = 144'h00d10286f5aa07330421f9db0422f5e8099d;
mem[61] = 144'h0ce70977fbeaef76f2fcfc7bf8bef63b020b;
mem[62] = 144'h0b1ef73301bf072ff4540718f5400049f59a;
mem[63] = 144'h109c0dc0f5400711fb6e03fe02190198fa50;
mem[64] = 144'h02120d77053dfef00d140d8ceee3fcb60c77;
mem[65] = 144'hffe2fd76f2330333f1b602690b1cf3abf501;
mem[66] = 144'h033008820be8f049efb3031ef81dfcd5005c;
mem[67] = 144'h010b0d32027d050ffffa019c0e4c0fd30d6b;
mem[68] = 144'h0b440fc4f35df66ff9850ad9f5caf7860265;
mem[69] = 144'hf71e03a7031b01630dbef619f2cc0d1903bd;
mem[70] = 144'h075a0d79fe0203eef4620eadfcb6f691f223;
mem[71] = 144'hfab4fa1aff6afbb5f72201f8f044f4640eda;
mem[72] = 144'hf665052b05e4f5c4f9dd013b021c048e06ae;
mem[73] = 144'hff2ffabeeff2f12bf506fadef755ff79faa6;
mem[74] = 144'hfb8d0bbc0200ffbff659f129f8370d770a83;
mem[75] = 144'h059a0b5ef10ef9c2fc3df475f1a70027f2a1;
mem[76] = 144'hf2e3fde9f147f718fa9af064f2e10ca6fd44;
mem[77] = 144'hfb690e3df456fcd209e4fc6c084302d7f783;
mem[78] = 144'hf672069ef39d0e27f317faac01f60c450bf9;
mem[79] = 144'hf0a00e2f0f24fbf2f60e020d02080cd3f8c1;
mem[80] = 144'h0bdd0cc40d410c67086504e30bbcf167f588;
mem[81] = 144'h09cf002409fdfcdb0970f125f479f65306a3;
mem[82] = 144'h0eb8f20708d10e17fab8072d09c10e4affaf;
mem[83] = 144'hf749fc48f8fb076af7cd09f3fb2ff0a803d1;
mem[84] = 144'hf22a0b09ff54fd1007c509e10b0af856f330;
mem[85] = 144'h0a6307cc097303b70b27fde70d09fe1ffecf;
mem[86] = 144'h022f0273076f007a051407330d77f04005f2;
mem[87] = 144'h0a76f695ff33f7820f9504810c180b73f4aa;
mem[88] = 144'h0d17f7230e760bfb0aee05a9071af0470e34;
mem[89] = 144'hfc99036506610abef9620583faa1fd5bfeac;
mem[90] = 144'hf257f224f0fe0315f8cef9f5f198f957ff79;
mem[91] = 144'h0e3bf7b70741f5e2f9defd0bf10efab3f586;
mem[92] = 144'h05950dfaf4370d69ffa9f8d90f43fb75f1ec;
mem[93] = 144'hf88d0d2dfdd2f357f856ff5802a5ff7dffc2;
mem[94] = 144'hf15afbad079a06300d35057ef0b8f6770468;
mem[95] = 144'h0ee2f4d502740a4002b0fbf503b2f23ef489;
mem[96] = 144'hf8a40fb3fc4c0988f5a6f630feb006aa0927;
mem[97] = 144'h0f76022cfa3902b104f4fa0a0cdd018df002;
mem[98] = 144'hfbaafa35f5fff253f271fc6304cef910f62e;
mem[99] = 144'h0e36f547fbc20141031e082c0921095ef434;
mem[100] = 144'hfd0dfd52f6810a0309e80a27053c0f4af179;
mem[101] = 144'h087b0c1af986f126f604f1c6059f09c30892;
mem[102] = 144'h05f3f0b301ddfde6faebfa1a06bbf26cfaac;
mem[103] = 144'hf12f01c80017f190fa910c690cb0f3690da8;
mem[104] = 144'hf97ef85ef08e0f390c2ff482fd49f4d009cd;
mem[105] = 144'h01800ada0317f8d7fe510f58f3e6f32ff316;
mem[106] = 144'h019df2fcf52309c801d6f70dffd5f4d30246;
mem[107] = 144'h0343faf401d00eac0be1071dfaee091d0793;
mem[108] = 144'h05a3f24a09dcfdcc02b70b76f51a012ffdb6;
mem[109] = 144'h02d70f260075f8930759fe7bf3dbffe20382;
mem[110] = 144'hf204fec2ef4504f80a85f892fae0fb70fe57;
mem[111] = 144'hf886081d01bffb4d00bcf8600118f619f959;
mem[112] = 144'h06bff253f96ff58defe1fc5b09c80816f5f1;
mem[113] = 144'hfabcfdf00305f01f08ce0ce4fd47f705f21d;
mem[114] = 144'h0b6cef7a0e13fc9ef5ad0e01fe600b7bf9b2;
mem[115] = 144'h05d701280a3df8c2ff42f79509e0ff050cde;
mem[116] = 144'h03be0e6c0d9a00dffbee033df2b00c0d063b;
mem[117] = 144'h03950469fed50b4af4caf2d30116008ff27e;
mem[118] = 144'h02d50adfff8d0c59051b0ab6fefff81df66d;
mem[119] = 144'hf006f1020b37fb340d7f0f1c0f3b0872f9e5;
mem[120] = 144'h0a9afae9efda0c00f49ffbdbf2db0721f920;
mem[121] = 144'hfc79f5b00bf4f1b7fba40685f5af0839ff39;
mem[122] = 144'hfbcc0e5e077402d9fbbe0a6cffd9f503ffdf;
mem[123] = 144'h0c1702d0f03bfb5e044302e8017309f9fca6;
mem[124] = 144'h0e300e4a028bf8c10d2df3c7f55bfb22fd00;
mem[125] = 144'hf88d0e94f5c807aaf7acff00f2bc06ed0d86;
mem[126] = 144'hf8cd01bb01ad0ca8fedcfdb10af6019ff79d;
mem[127] = 144'hfd4700fcfef70e2405ee0b9f06dbf8fff8a3;
mem[128] = 144'h07950bf40c58fc77f66902a80dfdf118f7c0;
mem[129] = 144'hf5b6faf50325f37f05020fbbf3a8075df449;
mem[130] = 144'hfe95f12c0997f7bc0230ff3b0c840a1704ed;
mem[131] = 144'hf822f6eefa7ff3f4f3a00a0ffc59fe9b0e90;
mem[132] = 144'hfcb7f97ff767f43c0b11fd3cf51b045d0c1e;
mem[133] = 144'hf74df2130aa9088dfe5903caf6d801d4f48c;
mem[134] = 144'h095e09a002f301bc00ccf3a004b307f305de;
mem[135] = 144'hf3d5f6effde4f5df0f1302040d97f5ef0f20;
mem[136] = 144'h0ad7f0db03f40af104e4033bfd2cf3330aba;
mem[137] = 144'hf3ad09e2043ffe3f02cb03b309110cc7fd79;
mem[138] = 144'hfac70576f05308ee065b004af8ecf92103af;
mem[139] = 144'h01b6f3e1fc28029af242fc3dfc4905def3e7;
mem[140] = 144'h057ff90c0269f916ff080140fcbdf26c09d6;
mem[141] = 144'h0175f830f82bffce0dfc0b1906f105d6f2a9;
mem[142] = 144'h0336ff58f7d20cb6fb580106fdd4f3adf2b0;
mem[143] = 144'hf74e002b0ddb08b001cafe0ff7510191febe;
mem[144] = 144'hf2fdf453018b0d2302bf03dcf3bff24103cc;
mem[145] = 144'hfa070f2904fdf0100ece032f05c6fbe4f6f1;
mem[146] = 144'h04cafcca0d84f4d50f67f5a30176021a074d;
mem[147] = 144'hfeb7016df1d6f499f46f07c7f128f4dd0b68;
mem[148] = 144'h090dfa1a0277f72b0a37fa2f00c6f0cc0b86;
mem[149] = 144'hf28f0a650f99ffd308fb0f8908960bd5f76c;
mem[150] = 144'hf703f0d60581efb9fd80f246ff53ff1a07fd;
mem[151] = 144'hf00ffcea0c86f5b209c8f0e80e63f4280ea7;
mem[152] = 144'hfb9402f8fd44faf104c5f26d0526f372fb2c;
mem[153] = 144'hf90c0f20040cf3f0f2d8f139035a0ce00673;
mem[154] = 144'hfec309310c69ff4c0b9dfb9af58ffe68f74e;
mem[155] = 144'h00ae0046f2c20d1b0b3a0ce805110f9f053b;
mem[156] = 144'hfd77f854027005bcf657fa51f1e4f69bf907;
mem[157] = 144'hfd9d0b790ef30183fe38018e0495f9fefbad;
mem[158] = 144'h04c1fbb8005409db0657ff65fa44f88c0350;
mem[159] = 144'h0490fe3b0d99f03af13afb8dfce50b630bd3;
mem[160] = 144'h04050a490398f8810298ffb4fe0ff62c097c;
mem[161] = 144'h0fbc031609c1f839028206befa0204ac0e00;
mem[162] = 144'hf66a0114000c0450f5a60c80fc6808abf652;
mem[163] = 144'hf7390becf49af257f67b08ef00ff01870e44;
mem[164] = 144'h0c15fdb20c55085afcd407fe0efbf42afc2a;
mem[165] = 144'h0ef3062408a8020c0e000129f5940b9ef812;
mem[166] = 144'hf2c10eab0e0e0afcf705061d0267f00e00fd;
mem[167] = 144'hf3ff047e01570834f70c0fb6f493fa06f630;
mem[168] = 144'hfa890a280cca0dd2f94b0a21f5ba00b40d52;
mem[169] = 144'hff86ef59fec40a41fb7408f20e8ef9380c70;
mem[170] = 144'h025bf63b01850657fe45fb49ffb0f81dfd48;
mem[171] = 144'h0932f7ee0b670dd90a64fef6efd00553f380;
mem[172] = 144'hf20c0bef09010ccb041502c0f217fe2ff9d8;
mem[173] = 144'h0474f9330981048c043c09d504e8fd320343;
mem[174] = 144'hf04702990839f14c0800f8bbf76df23efbb6;
mem[175] = 144'hf38bfdc9fd8207fffefcf0b00b840476fa53;
mem[176] = 144'h0e6dffb9fef6fdec03dd02e0fa75f833f38c;
mem[177] = 144'hf283086ff8fafe0bfcae01200754ffb0f5aa;
mem[178] = 144'heffe0d40053508be0bacf90103760497f0d0;
mem[179] = 144'hfdb407760f120b09f68c09feff35f869f0f9;
mem[180] = 144'h015b0d7cf528fb1707a3f4e8f07f0b9705e9;
mem[181] = 144'hfd0ef4ad0ed7f1ccf242f95cfcddf674f115;
mem[182] = 144'h0606f8c608b9014104b2f21ff811f83bf6d7;
mem[183] = 144'h0ee004faf9aa09affdd4fb34093303e9f54a;
mem[184] = 144'hf0b20aa2f9f4056e05ea0cef05b40f0bf35f;
mem[185] = 144'hfab408eef2cbfdd9f8af0676f423f853035a;
mem[186] = 144'hf4a4f882f276013308d3f460038ff712ef88;
mem[187] = 144'h08c5f26a029bf9fb08d80d990070fad5fa70;
mem[188] = 144'hf86bf95c045af2a30305033807b10850fe9e;
mem[189] = 144'hfa060044fcf803faf0dbf9e80be6f9090bdf;
mem[190] = 144'hff7ef43ef27d03550630f9d00a32fbac0952;
mem[191] = 144'hf92af59cf2f9fd160a12f646f8870332000a;
mem[192] = 144'hf1c706360643efe5f95207ff0b32f65b006a;
mem[193] = 144'hf2000c2e0090f1d8fcb2058f0b7af2e50b34;
mem[194] = 144'hfb07f418fdd801350acd0dfefd62f15e05a9;
mem[195] = 144'hfc930713f409f9300700f2a605660028088b;
mem[196] = 144'hf7640c2d083af9cb0a0d0d46f1730f39f3b6;
mem[197] = 144'h0ef90bdd096606e40c5bf11e02d3f3440ed3;
mem[198] = 144'hf7490af2f0a8f71df0320d8408b40b59f1f8;
mem[199] = 144'hff400751f3ef044dfdbf0876f49bf888014e;
mem[200] = 144'hf6befc0707820b6effe803d106f9f86001d7;
mem[201] = 144'h049ef3e5f27ff46a0b57f5080bf201ff0561;
mem[202] = 144'h0c0b0f0df84dfb9804410e04fa49f5df0983;
mem[203] = 144'hf79e0250fd26fe130680f0c70ef8f790ff15;
mem[204] = 144'hfb7df4e9fb240c4e02130fb90ecafcaff188;
mem[205] = 144'h0b6f09e8fe140827074a06c90c0e0477096f;
mem[206] = 144'h0db4f2840e0501d10e13034d0d1ef504f070;
mem[207] = 144'hf6affcd2f5d6f6090762fd4cfbb2fdd5fc0e;
mem[208] = 144'h0ae9f2def46af096fc42ff80f38f0bf9f5f9;
mem[209] = 144'h0aa600c9f566f05d0a100a090ee5f18f08e5;
mem[210] = 144'hf3d10374f12d0664fb8a0fc40b24fd5aff8a;
mem[211] = 144'h0741068ff8080a6f002603f4f66f0553fc80;
mem[212] = 144'h04c80299fbb00b300dd107280b21f09b0724;
mem[213] = 144'h02100e81fbce019a02400f780a1dffe0f22a;
mem[214] = 144'heffe082cf0f8fa73f2fa0863f4a20e56fc56;
mem[215] = 144'hf4e2fcab004c03a501be06d8007900840d85;
mem[216] = 144'h06ff01e9fe46f708008109f0f36604e1f794;
mem[217] = 144'h02b80d69f0f003defabb0fdbf666f354f715;
mem[218] = 144'hf693ef1bf5c2045bf778f582f1370399fb1e;
mem[219] = 144'h0b450d1d0bbc033bfe4e073d0cccfcd60dc5;
mem[220] = 144'hff4e0d630e730ba3f631015cfe24f715f74c;
mem[221] = 144'hf6b4002009260b0a0803f578fdf008a10347;
mem[222] = 144'hf35c0ce7fc04f7320ac309b3ff5efe730c5c;
mem[223] = 144'h037df66ff91f055f0ad0f54109e1f356f23b;
mem[224] = 144'hf961f420087a0bf8fd61fe850bcffb0b0a9b;
mem[225] = 144'h0255f9bf0b1c0419f340f9ae0cbff4940753;
mem[226] = 144'h09430032ffd4eee4f145073ef9cc0eb7fa2a;
mem[227] = 144'hfc39fd2df7dfff650bce013ff4050e3af8d4;
mem[228] = 144'h0ba302f5f71f03aff042fcd7f8770ecd01d0;
mem[229] = 144'h02a0fa1408420e8909f4fabe04a70e5af942;
mem[230] = 144'h0287fb5d0c830c420dd10d4b0465097bf3c6;
mem[231] = 144'hf6ccf2c1f3ddf85a04bbf9480121f992efa8;
mem[232] = 144'h0c3defbbf3cff0cefa3ef8e7fd5d094c0c95;
mem[233] = 144'h0c9008dbf3f709cefe64f9ccf5c0f68d0c89;
mem[234] = 144'hf0f9056df5caf9b901800a5a09acf85df56b;
mem[235] = 144'hef89fca7fbf0fc9604b3f71c0e2d02b2f843;
mem[236] = 144'h0db80662ef32f1b9032aef9ef1eb0a9e0590;
mem[237] = 144'hf72bf2fff83bfdad031a060802820318f93b;
mem[238] = 144'hf083004602360042f2e2fc8fffe40bcef252;
mem[239] = 144'hfb1df748f204f4fcf29cfdbf0c9e024ef0fe;
mem[240] = 144'h0d50ffe7f57c0616f9c10a79f8ee078a0335;
mem[241] = 144'h05660e49f4770aecf4d50ef2f501f02df74b;
mem[242] = 144'hfd7b0c33038bfd6e0fc6f23bfcf3f032f733;
mem[243] = 144'hf014f873fa1af1860c83f9abfd9609940062;
mem[244] = 144'hfb27023dfb790063fd12f1dcfb76f2d40ebc;
mem[245] = 144'hf1aefdc5fd75f12e0e6207b3fb01f7b9fd6e;
mem[246] = 144'hfaa7048ff1a0f2b807cf0db6fa4df6c8fbd6;
mem[247] = 144'hf79d0f150d4bf3d3f5f80c0e0f5cf75ffebf;
mem[248] = 144'h005707ac0443f761f151f00902c50eb30225;
mem[249] = 144'h0b9cf6cf01440117f2b1f47500880b3e0962;
mem[250] = 144'hf87ffe00f031040bfd7b0f55fa950382f78e;
mem[251] = 144'hf4f1fac5003cfbb10dcf021e00bbf6fcf00e;
mem[252] = 144'hf4ad0be20c29f0c500080a4a020f0a6bf70f;
mem[253] = 144'hf10efc9809b7f313f3e9fe16f75efede0cc3;
mem[254] = 144'hf1b9f73408e30dca044405e5fad5f5c009ff;
mem[255] = 144'h0d3df166f9aa0e80f7970585f73bf40af08c;
mem[256] = 144'h00a5f37d080bf690f90efdc3f680fb230c0c;
mem[257] = 144'hf074f91706eaf5670a65f320fcedfae70262;
mem[258] = 144'hffd60e82f433fbcbf9fe03a9f3640783f439;
mem[259] = 144'h0f06f8760b0607fe0e49fa7d01d6fff3f6d3;
mem[260] = 144'hf5e8020308c3f7d606b2fc0c02bffdbafe26;
mem[261] = 144'hf7f5044e0322fba5fac4f29efcde0cf5fe19;
mem[262] = 144'hf28ef181fade06a9f4f00a97f78af2b8fd12;
mem[263] = 144'hf1df04f5f43cf4b0f074f2c9f69b0d1dfc26;
mem[264] = 144'h0c3ffc9f067b0ae6f7a40dfaf22f08ebf485;
mem[265] = 144'hf665f1acf5caf3c205a3f3a30d3e0d6dfd07;
mem[266] = 144'h0356075b051c09340a3b0aebf83700a80ab7;
mem[267] = 144'h0e3a07020472f0f8fca306a903b3f940053e;
mem[268] = 144'hfc0bf7d40b1c0422f5faf0150ddff1560241;
mem[269] = 144'h0841019ff9d6f8c1063a098ff0fefdbe0a90;
mem[270] = 144'hf7e9f57cf624fc240c53f6a3f34f091b0040;
mem[271] = 144'hf9970d7d0c38fe000d73fc7d0efdfba6fc3e;
mem[272] = 144'h01acfa4dfc000486efb406d7024df60d0e85;
mem[273] = 144'h0de700c507b0f9b809ef0218fb20ffbb0767;
mem[274] = 144'h07daf3e8f073f498f020f161f61f077e026a;
mem[275] = 144'hf267001c0fa7031efa1004660142f6f7f353;
mem[276] = 144'hfa2609c1fa3c08250a010aa30250fae00909;
mem[277] = 144'h0975022cfdabf18ef8df04adfd86073800e0;
mem[278] = 144'h007afa40003ef15a0f38f3f10ded023a0d24;
mem[279] = 144'hf58a06d408fa03dc0583f914f67e00baf49e;
mem[280] = 144'h027e08edfdeaf599fc6906d20547044df1f1;
mem[281] = 144'hf80f0a43f6bf0bc902b50d56f9280282fe5c;
mem[282] = 144'hef48f0a10b0704f7f22f08870416feedfe18;
mem[283] = 144'hfaa10756065401daf48efad9f5190cfaf6c3;
mem[284] = 144'hf74802dafab001eaf1c4fe66044dfe42fbba;
mem[285] = 144'h0ae008ce0c3c063306920de4fd62fcd60d4e;
mem[286] = 144'h02c2075e029d0c9000c60c3e0ef7f5aff25a;
mem[287] = 144'h08b30f3df16dfc360cdff7b60ce4086c075e;
mem[288] = 144'hfe9c0b8dfe6df442f648f8faf292fd4109cd;
mem[289] = 144'hf37f0ac3f42105bd06e1f65cf242f053f8e8;
mem[290] = 144'h08910666f53a0cf1f2c8eff10c7cf584f9eb;
mem[291] = 144'h0f5aff3b0ac205f0057bf7b0f034f90ef7d9;
mem[292] = 144'hfd6af160ffab020af37a0752f4defdd90824;
mem[293] = 144'hf55ff47b0da3fbe30c830e42f406f8f50965;
mem[294] = 144'hf739042c09ed0a2c0cba01e5015b055efab5;
mem[295] = 144'h0b10fad104bd044af209010f038efc19f9ca;
mem[296] = 144'h0815fcd4f550ef88f7e9ffc5efed0b78f8d3;
mem[297] = 144'hf766ffcf0b7d0405fd890151f5530833f375;
mem[298] = 144'h0d28f9f8fb2b061f06def882038bf5680122;
mem[299] = 144'hf05bf6d6fbecf3a603bcf0aaf3c80235ef90;
mem[300] = 144'h02bfff5902cdfd76f4f4f302ffddf3d707d7;
mem[301] = 144'hf7fd075feee5073701bbefbafb2af091fcbe;
mem[302] = 144'hfff4fce9fd0a0b1801daf57f0150f62c096a;
mem[303] = 144'h05650e2dfe5ef6acfd1203c900ab0a32f742;
mem[304] = 144'hf7d2ff38f6080cee04eb09630efef434fa75;
mem[305] = 144'hfac6ff3b027df2360bd20a9ff27ff487fa86;
mem[306] = 144'h03a2f76ff2c10a0d08f007940472fd0ffa4f;
mem[307] = 144'h0f8e001005fefed90725f3a20c500997fdb7;
mem[308] = 144'h071d0d79f272f5230655fd94008403440768;
mem[309] = 144'hfb32fd4cf47b0fb50c710745fe8007800c02;
mem[310] = 144'hf6f7f512f3a5fd01073d054ffba60548f3b2;
mem[311] = 144'hfb17efd5f97ef79e008bfaf8050c08850bca;
mem[312] = 144'h06a20a2bf35805aaf28d0d20fd7bff67f402;
mem[313] = 144'hf3b6f1d9f7f105fe097107d0ffb3fa3df8ad;
mem[314] = 144'h0bfd0e06097e09f1f81af4ef05a2f88a0a04;
mem[315] = 144'hf16ef5d60980f3530461012af465f6ae068e;
mem[316] = 144'h0944fb960bfa0dcff5be0eb301820ed90470;
mem[317] = 144'h06800124fcbd03cc03ddfab20a1707ae0c91;
mem[318] = 144'h08b50806fcbd0f670c49f98df465ffddfd7e;
mem[319] = 144'hffd402c60556f4c4f642076cf38ef5bbfad4;
mem[320] = 144'hfda30a93089bff7ffde0055af10ef215f594;
mem[321] = 144'hf356f455f24b07770caff2bd07fb0b9ef61c;
mem[322] = 144'hffcaefa8f756f3c00b28f257fcab002cf85f;
mem[323] = 144'hf5dd028b0ea701a00198f7910ef9f14d018f;
mem[324] = 144'h0e040a62fcfe0957ffb30241f543f58bf684;
mem[325] = 144'hfb61fb4bf72503c90b1dff1b0633feb80875;
mem[326] = 144'hf23afc2af2850987ff6a0724f065ee5af0dd;
mem[327] = 144'h0193fec1ef98030afc410be2032a003bffc4;
mem[328] = 144'hf24af89b0e9df21907b3f66d060a0abafcb3;
mem[329] = 144'hf585f9290140051809080eeff92af7b5f96b;
mem[330] = 144'hf2510eac0460f8130af1f1edf2d3f6e50b6e;
mem[331] = 144'hff2e0b2df617fb2107f805be01a6f0b1f741;
mem[332] = 144'hf91f02f3fecf06730cd4ef72f056f3ee0cd6;
mem[333] = 144'h0e6904d009c90353005103210476f81bfeea;
mem[334] = 144'hf7680363f190f3be0708f178fa2affe5fb04;
mem[335] = 144'h0749ffecff08f4220e4a0427fe8b0e3702bc;
mem[336] = 144'hf94909f7f61ef6310e650e2308ab010aefc1;
mem[337] = 144'h003c0dcff103080900750142ff69f5c5f510;
mem[338] = 144'h08de04e3015901eef094fa610c11f69af9b0;
mem[339] = 144'h0aa5ffc908c604e80f7f01a5088efd3bfc14;
mem[340] = 144'hf146f510f5d60a9df45af790f02cf607f09e;
mem[341] = 144'hfda504630d9500280e27f2d4fd920785fc6b;
mem[342] = 144'hfc02f109f205fe6dfb46003d06650755f48b;
mem[343] = 144'h0150f6830789f5baf4cdf0f4f8420fa7f189;
mem[344] = 144'hfa2c0038070d04d1ffd2fe830bf60ceaef0e;
mem[345] = 144'hef150be907ea0c59efe20e63fa1f0088fcde;
mem[346] = 144'hf101f28d09ce0f3b08550a5a07b3fc92f252;
mem[347] = 144'hf62801b2f85f0bce09620bfef6a007390772;
mem[348] = 144'hf87902dbf642093ff44ff3dbfb1a0b08fe71;
mem[349] = 144'hf735f8b6f6cd03acf885fb76fc36fe210a3c;
mem[350] = 144'hef13fc100e67f7ba00adfad9f2090c27fe4d;
mem[351] = 144'hfe2d0b3f0448fea3f63d038b080bf2dcfece;
mem[352] = 144'hfeeef93c07b8f9ebff70046c0ed70437039f;
mem[353] = 144'h077109e70ac6f351f652035b0d77f4ad0264;
mem[354] = 144'h05e6f5d1f64c0596f5400d2605670adff0d8;
mem[355] = 144'h000df689f014f65402a5f8a0006af70a083e;
mem[356] = 144'h0d6bf2a00daaf95c0bddf6f20b730f81f659;
mem[357] = 144'h017801a40b570651fbb5f5d9f4f70fa108cd;
mem[358] = 144'hf2c00e89fc03f342040af698f28600baf471;
mem[359] = 144'h0d1c0c69ff3bf00e0f0bfca40b94f82b0b5a;
mem[360] = 144'hf9d20e6f0dc6f218fba6ff84f29401110e77;
mem[361] = 144'hfcc6f698f2f0f0910e0b02ab0b96fc390581;
mem[362] = 144'h024ef7d507a50144f8900e6d03bbff9f0a1e;
mem[363] = 144'h091604c2f84cfce9f6880ad2efbf0b5a0e54;
mem[364] = 144'h02770c360576f5550613ffc80050f78703a7;
mem[365] = 144'h0e21ffce0c5e07b90523fda7fd7301730d47;
mem[366] = 144'h092cfcccf673fc2bfad50448047d0941ff39;
mem[367] = 144'h0e8df258fc27f849f1d40c5309fcfa1c0961;
mem[368] = 144'h004d0ddff90c023e062f06dc0778f64a01db;
mem[369] = 144'hf79205910bb90a0f00c8f6ac01500d9e032e;
mem[370] = 144'hfe50f35e0f52f28b05de00c1f1dd027df202;
mem[371] = 144'h0dfb0c8a0051066d0c29f35ef8f906a507d0;
mem[372] = 144'h037ef55df1b9068cfbe1f4a000be0445f1ee;
mem[373] = 144'hfbba0a30022df977f6e5f8f20cf7fc430cca;
mem[374] = 144'h0b52fef10c8c0491f803ff2b081ff4730811;
mem[375] = 144'hffbdf251f97a084b0d6bf02a01f50bdd0251;
mem[376] = 144'h021aeff40d020e72f85cf6ed0abff3370319;
mem[377] = 144'h0bd402b80ac6f85a094ffad8f5a2f81ff323;
mem[378] = 144'hfa0cf184f33ff6380867fdcc09fff8180c89;
mem[379] = 144'h0f82018d016af623073a011d0d4af6910abe;
mem[380] = 144'h0eaf06a5f7fc012002460c37f74b0365f40e;
mem[381] = 144'h09e30150fc06fa1eff4e044c0e95fdcc0289;
mem[382] = 144'h0f53f37f0f76f66ff19c08c4f7a6f951fdda;
mem[383] = 144'h0154fa98ff5b06cbfc9cf627f3b2f8410d2f;
mem[384] = 144'hf8a00834f5290678faff0b9d0e04fa4e0e6f;
mem[385] = 144'hfd23f4fd02deffe7fe8f061101f9fcc1fed2;
mem[386] = 144'h0c2feffcf63ff6f1f1ba09d003a3f000fedd;
mem[387] = 144'hffac0c56fa1b0b45fed0f834feb1015cfa43;
mem[388] = 144'hf25bf3eaf4b5016e0b20fc30fb7b01f0096e;
mem[389] = 144'h03dff0a007c3fa910c01f1720005f09cfb74;
mem[390] = 144'h0763f8e2f903f720068af7bbf2fa0505f1fc;
mem[391] = 144'h017f0596f4370e4300a40f9ef6da0d96fb9d;
mem[392] = 144'h0e23f4b1f63400acfd980135f8c4091302cc;
mem[393] = 144'h0a6d05810481fb12fe80fe9c0dc6fc97fd59;
mem[394] = 144'h0ed40f3f02c2efbafa50fc140f490f81f3bf;
mem[395] = 144'hfd6dfee609fd0875f41efa4b03f5fa680db3;
mem[396] = 144'heff00b4cf255f46cffca02f6f4cef6f70696;
mem[397] = 144'hfba9f6b809ab0216fd8701d30c840d4c018e;
mem[398] = 144'hf9d005e00863f2ac00cffde60ba308d0072f;
mem[399] = 144'hf47809d30bc0f04ef7e7f3050f40028f0db4;
mem[400] = 144'hfb3e0422fb6aff8402b704a3ff6d037d013c;
mem[401] = 144'hf88700610b9ef2acf40ff2f2f4dbfb6e0c48;
mem[402] = 144'hf13bf6a90b5202ebf38e02eef43f00b4f55f;
mem[403] = 144'h090504d4f9e40f41f829fd7ef4a503a8f36d;
mem[404] = 144'hf99bf4f8f04301870a9b09df0f7f0d5c032f;
mem[405] = 144'h0e0f0613f2600c2ff90c0854f07ff1500567;
mem[406] = 144'h058b0ab000350c56f3350e97fed40777fbc0;
mem[407] = 144'h0cb1f3f2f7d603e200bc032301c60b3af054;
mem[408] = 144'h008df78ff401068c08e90652f258f547f91d;
mem[409] = 144'hf42909b600d2f7af0f380781025f013b0f42;
mem[410] = 144'hfbc8f6c6ff130f04fca70e01f1340f62f31d;
mem[411] = 144'h02c9f8a40cecfe7a0563f31bf3fef888f87d;
mem[412] = 144'h0d91f2bef26bfc1e0dc80548f41403240528;
mem[413] = 144'hf00afe270a2602140e8bf035f9f7f6b10467;
mem[414] = 144'hf0bc0353fa51fdd4f1880ba60f5afd91fba2;
mem[415] = 144'h04f9f7b6094ffed7fb1fefe9f331fda8f83d;
mem[416] = 144'h0a29f586f824075ef40dfbd6070c0487f5eb;
mem[417] = 144'hf447f706fe7a0cb9f4acf0d608d4f5e7fda0;
mem[418] = 144'h00d60546f731f105f7bdf139fd5a0dec0a92;
mem[419] = 144'h02140e1e0d70012707e103b8fe5ff547fde9;
mem[420] = 144'h0ea10574fc880fd3f2d4f3b00fed083e0c5d;
mem[421] = 144'h04c70aec0e430590fcb10697047f02b5f431;
mem[422] = 144'hf3fef74d09c9f6770d8b0c20f3b7f29bf1e9;
mem[423] = 144'h03d0f205f3820269fe420e570b83f868f41d;
mem[424] = 144'h0f30f25d0a5df1e7055401e5fd64f730fb0d;
mem[425] = 144'hfa5502f3f91503f3f8ddfb2e06f90a01f9ba;
mem[426] = 144'hf202f4c7050c0b8d0f5903970c43f103f82b;
mem[427] = 144'hf51af3fc0ebd0d8ef2b00f3ff36200e90813;
mem[428] = 144'hf92b0e550dc0032b0003f09a0dfb05effbf7;
mem[429] = 144'hfe95f636f7c40109fd0809f105bd01770ab0;
mem[430] = 144'hf13b0dbafe8707b80cf50308fe63fe070339;
mem[431] = 144'hff2cf7a10f03019af7ae01410529f805fc3b;
mem[432] = 144'hfdd3fc18015d0c17fa9309e20fb1ff57f2b1;
mem[433] = 144'h030af8bc0fa601d4f70ff031016dfdc50ccf;
mem[434] = 144'hf4b0093e05530bc405fdf73ffbb105ff0a01;
mem[435] = 144'h0394f54809b6f8fcf01700b00e7c0ab309d3;
mem[436] = 144'h0de5f01a0554faf0064e00070e5403ebf18f;
mem[437] = 144'hf689fb3605e90f21f556fa2c0c8efbc9fca1;
mem[438] = 144'hf736f8520df4fca209bef992fc85f5530a26;
mem[439] = 144'hf79001c7f8f7fdb8fbfdfb91fb96fc10fa29;
mem[440] = 144'h0db40192ef17effc0f48090af4a7f41c017c;
mem[441] = 144'hf9adf82feeda05d3fa8400c10afcf451fb88;
mem[442] = 144'h087cf0980c850a79fec9fd1f07b602080d3e;
mem[443] = 144'h03c1f5c2072c05c9f21b0779f7c70744fdd7;
mem[444] = 144'h081300170a74fa4bf833f298fce6fb0dfb85;
mem[445] = 144'h0fca05d604b50a50057f01730f5df88cfbe5;
mem[446] = 144'hf2090ca70d15f76f0d6cf71c0637f23a0c91;
mem[447] = 144'hfa3a088fefdcf6410613f1c40778fce5044f;
mem[448] = 144'hf65c0d85f30efac000e9f7a309db0f780b10;
mem[449] = 144'h0c080367fecf02d30a6afb6908e60d7c0971;
mem[450] = 144'hf7f2f9ce082f09a707b0fcdef98df40a0abc;
mem[451] = 144'h0154efc0f9db0685f3ef02780ebaf6adfe77;
mem[452] = 144'h0f350987001f088a06af0bcb0a190d3df11b;
mem[453] = 144'h07f4f242f050076a09b405bd0b880efbf3f0;
mem[454] = 144'h0f89f9f3ff2602d5061b0dd2fa5e03400e9d;
mem[455] = 144'hfe0b0ec700fe0802f78efc10f4780ce4f808;
mem[456] = 144'h06bf0a1d0f94fbf703ecf528fce7f132fb0c;
mem[457] = 144'h030400dbf750018ff902f4e10e6e09e40833;
mem[458] = 144'hf3ae025704f402b20bb50ac1022507b90f0d;
mem[459] = 144'h046f07fcf25e0d06ff5efd03f262f760f3fc;
mem[460] = 144'hf0110a44075afca10141fa11f85cfb19f47e;
mem[461] = 144'h079d0cdc0e98f2f90a2b088c02640ec100e1;
mem[462] = 144'hf267ffccf360f698f41e0d80f8b4f993f948;
mem[463] = 144'hf5a5f2890115f1a80c40044c0bd00f6607c9;
mem[464] = 144'h0273066a0bc6f63af503ff6408a30455f489;
mem[465] = 144'h07a60736fa81f779f5d2fd6f07eff62ef6f3;
mem[466] = 144'h0238f22604150e97f553097bf772f4dd08fc;
mem[467] = 144'hf64efa1df4c9f7980f20f2d40a83f38709fb;
mem[468] = 144'hf69dfb11f49105a8f9fe01e70ebc0bedfb4b;
mem[469] = 144'h0cc90e770de6f714f80efde0f32e00c0ffa4;
mem[470] = 144'h08200514f9e401e705b5f6c7046df8d6fd38;
mem[471] = 144'hf88bf6c10cde06aef3ce032bf770f30d007c;
mem[472] = 144'hf79a0a9e017efbd603a2f4330a98fc16f895;
mem[473] = 144'h08bff873009bf1cdf4ce011ffe670715f43d;
mem[474] = 144'hfb73f7b0024cf85d0401f605efdbfd58f48e;
mem[475] = 144'hf8d308910ddb08c1fb1bf7aaff41ffd6059b;
mem[476] = 144'hffb6f7aaf1a4fd48fc0e09fc0afaf67a0fcd;
mem[477] = 144'h0d5008ddf5200a8502e9f5ebf182fc05f8db;
mem[478] = 144'h04ccf9ccf58001b1f3780de2f6c9f091f525;
mem[479] = 144'h0ebc0cbff3e90c5a0eeaf6e5f782f3b5efaa;
mem[480] = 144'h08aaf4faf31c0946fddb0844ffb9f8f9f53e;
mem[481] = 144'hf9c3ff080c73ff99f6c20e2408880839f284;
mem[482] = 144'h0b77f3dcf956065ef7e0f81e05f4f36cf7dc;
mem[483] = 144'h031ff287f8770a59f6b70723f340043ef135;
mem[484] = 144'h0ea9f6eaf5aa02de08b5f397fc920c92f3a5;
mem[485] = 144'h0e45ff6504ed087d04c9fd8f0f3709300632;
mem[486] = 144'h0f86ff77f0b4ff83f7f6f3350d4ff697f383;
mem[487] = 144'h022efc0efca4f0f5fcabf10d05b80aea0a2a;
mem[488] = 144'hfe700b0f09a4f074026c000f06e1013c049f;
mem[489] = 144'hf7beff07f34bf13b08ba0d58fd2b0158f423;
mem[490] = 144'h0a1d0d0cf8d4f81df6530ba1ff5efdacfce4;
mem[491] = 144'hfc3dfeacf2a4fb020c6efeb205620727f6b7;
mem[492] = 144'hf0c1f6100752f22202b70828faa5f5dcfdbd;
mem[493] = 144'hfca9f0020f3aff94f1ed0c21f1350f9df13a;
mem[494] = 144'h0c6601d2f3af0272006c0b250e0df1d9fb36;
mem[495] = 144'hfd27fdbdf603fcf60aaeff08fb18048dfe8c;
mem[496] = 144'hfa420934fe53f06bf4f0f3bff76603eefb0a;
mem[497] = 144'hf323f66a0182f0340baff9def68a0467fc30;
mem[498] = 144'h01e0ef22099c00ed061c074efc6a01df03e8;
mem[499] = 144'hf2b0f858f482f957024cf48af8940454ff23;
mem[500] = 144'h0d140652fb35f873f92600cbf048f219fc32;
mem[501] = 144'h0cbc0c48f6390465f855f278027508a9ffd2;
mem[502] = 144'h04cc09b1f25ef3f8f563f1e80668fb5ceff6;
mem[503] = 144'hf984fe56f151f0be03490f1df0d805d800f9;
mem[504] = 144'hf40bf74502c00da60ca60942f8c7012d095c;
mem[505] = 144'h050ff44ff9890a770edd05940e250565031c;
mem[506] = 144'h0540fb1c0c070e5c03a5f6c30277f6d509d0;
mem[507] = 144'h00b10477fc24f6f5fbdd052f0b1efbecfd46;
mem[508] = 144'h0206ee70ff220be9fd1ff43403cd020407b1;
mem[509] = 144'hef90f28dfaca07e303860e4a0264f5da0dae;
mem[510] = 144'hfb0ff0f20bfffd34035df46a01cd0bcf09d6;
mem[511] = 144'h02800ce2f9a8fb39f4cbfeb706780c73f933;
mem[512] = 144'h063b07e7f3bb01a6f64109b30773f976f845;
mem[513] = 144'hf041f0b5f26ff34a09ccfd61013ff79dfb85;
mem[514] = 144'hf2f30d7a0971fafb0e92f454fc7b02c10870;
mem[515] = 144'h0d77041bf3effcfef128f441f441fb04096a;
mem[516] = 144'hfbaafef30e12f4bb00b0083aff410d8dffaa;
mem[517] = 144'hf80ff508f5b509e7fa24fde4f253f7a9f79d;
mem[518] = 144'hf291f51cfbfefaa2fc080153f8ebf0400eb7;
mem[519] = 144'h0ea30c6bf32302c0033ef6e0092f02a600b2;
mem[520] = 144'hf7720bd7fd820a82f91ff640f45ff505fbec;
mem[521] = 144'hff75fd40f3b0f88ff0ef05af0ec60a03fdb8;
mem[522] = 144'hf85bfaea03820113efa80603f1b708b30514;
mem[523] = 144'h0944fd72070204e2fc9e0b37fd6d0ee108a7;
mem[524] = 144'h05730c14fe29f65df8c90827f413f9ab02e9;
mem[525] = 144'hf646f42b03d305e2f280ffb60d03071d0295;
mem[526] = 144'h0fa7f1aef269fd2efa80fcbf03690127fad9;
mem[527] = 144'hf977fbe0f7d00107fd42087ff2770c00f2a7;
mem[528] = 144'hf462f726fe4bf94802f50d2eff0bfeaefdc3;
mem[529] = 144'h00990c1c0210fd7702630668f48af311f231;
mem[530] = 144'h06630a28f2f3f28b09a10f03f74c04370a5e;
mem[531] = 144'h07f3fa490af8f63f04e1f989f7f60981f6ba;
mem[532] = 144'h031406b0fb0a0c72fad5fffa070c021d0a4c;
mem[533] = 144'h0d5ff103fe9ef65a0de1f8a20e9dfe830120;
mem[534] = 144'hf8ce04f6f572f8a50de0fc42f6000885f997;
mem[535] = 144'hf12befe4f3b2f8ba04a5fc68fc34fa5c09cb;
mem[536] = 144'h0e5d0e3008e3f57608db0135f299f4d6fa7b;
mem[537] = 144'h0b130b0af10704e1ff310906f2550e23004a;
mem[538] = 144'h063feffe06acfda2f1ddf9940e4a00650560;
mem[539] = 144'h0a15fa20fe500e980f19fc9dfb270d210233;
mem[540] = 144'hf722fe8afa71fa7ff9a10150f561f2d9fe80;
mem[541] = 144'h041cf44f0b04038006a8f7a9fe9104370b6f;
mem[542] = 144'hf9220666f957f1c50c8209effc49f6c6038b;
mem[543] = 144'hefbaf98ff49803d1f4d4efbeff20f9bdf173;
mem[544] = 144'hf64d000407f105a1eff7fe1af29df9a6f10d;
mem[545] = 144'hf0780416fd13fce3f33c027b06f803e4f26f;
mem[546] = 144'h05b0019f0a11f561fdbff0f3f6cffcc1f3e1;
mem[547] = 144'h0bb40c44f7a8f16907e1f1320530f450fe38;
mem[548] = 144'hf1480d2b0895f9c50b660e4205b30381071b;
mem[549] = 144'hfb7df7d40457f4ecf1d2ff050ca800160797;
mem[550] = 144'h0bf60688018303f3f76507e7f20c057d0535;
mem[551] = 144'hff11f954081f0b260a8d0550fefc020cfff4;
mem[552] = 144'hfb090ae3ff5905a8fb8508420a1b08f2f56f;
mem[553] = 144'h0c6b08e30c76ef28f20ef6700a980c80fba1;
mem[554] = 144'h0b43f93ff9cdf5bf0ce40e6300b60e120668;
mem[555] = 144'h0e340614000506f3052af34bff89f6c3f283;
mem[556] = 144'hf981f2e70ef8f0a3fd30f07df17f03140827;
mem[557] = 144'h0bf50f4cfa8bf5c00e320ca9f5c5053b0c22;
mem[558] = 144'hfa65fa85f5b0fe6e002401bef48c0dfc05db;
mem[559] = 144'hf5c3f948f18304e0fdbffcb107e8fcc8fe68;
mem[560] = 144'h045d071bf2d2062af0020eef0a7bf7a20059;
mem[561] = 144'h06f60a860fd1f5270de906c7f703fd3df5ac;
mem[562] = 144'hf396fad9007bfd8f095102d500520ba700ce;
mem[563] = 144'h0cc106930737f2d3f774fb16f02806ddfb4c;
mem[564] = 144'hf0de0bd00491fe1206fb01ac03d4f5b9f5b7;
mem[565] = 144'hfaa1fec6f61b0b7506320797f9a301d901e1;
mem[566] = 144'h060c0e70f6ee00cbf378fc7cf841019a08f1;
mem[567] = 144'h043f000a054efe39fda1f0ca0b53fc2cf0d2;
mem[568] = 144'h08a50016f04fffd708e3f4a1fb95f4e2f3c4;
mem[569] = 144'h0872fd00fc49f58df860f8f9f96c0cf5fe6e;
mem[570] = 144'hf11f09aaffa8fc95fc62fe1d07cffdc30cf6;
mem[571] = 144'hf21af5450687f9b4f7a3f5d5fa46fc44067f;
mem[572] = 144'hf5890ddb05bbf95006b602200158f11d0c2d;
mem[573] = 144'h0cb803700c660ae40fcc0bc7f5520694fa71;
mem[574] = 144'hf2fb02270101f3ebfabafb95ffab0d54f001;
mem[575] = 144'h05f8f2dc06d703a40723fe5a01a402cd0520;
mem[576] = 144'h0f4d03d5f7650749f0d9f2de0af2f882f397;
mem[577] = 144'hf22803c703d8097ff0edfb37097bf4d2f3e5;
mem[578] = 144'h0443fbef0c490b5a0a13fb3bf1460168087f;
mem[579] = 144'hf477f0cbf478f428fe3c0ea20253f1b2097d;
mem[580] = 144'h03eb0257f881feabefedf03b0c19ff870d13;
mem[581] = 144'hf6a60a33f6490789016d0eb8016e00d40a69;
mem[582] = 144'h034c095df35901f90e1e09700a36fbd1f213;
mem[583] = 144'h0144f891fb29057efdb507d2f2f7fb8efc16;
mem[584] = 144'hf068fd87f3bcfb22fdbefe2c01710ebaffb7;
mem[585] = 144'hf5dff5dcf68f09570e7c05860df8f93df12b;
mem[586] = 144'hf436fe68034f0450f2e70b2208950d87f9df;
mem[587] = 144'h0b22f105067403030dd6029907efefddfe6b;
mem[588] = 144'hf436f2a8f62df82cf665f9c20d4bf960f19d;
mem[589] = 144'h05b103fe0f1af5be0b37f05b05e6ff28fb0b;
mem[590] = 144'h036808a30364fa44fada0ac7fdd90e0c067c;
mem[591] = 144'hfa3d0130086e04e70cf5f0c60c1bf487f95c;
mem[592] = 144'h02abfc8c0d30f5760dea09ae058cff7befe1;
mem[593] = 144'hfb26f6dd03280c6af5490ca6fa0a02c2f042;
mem[594] = 144'hfcf30939fe810dfd03960595f489fb1e0e82;
mem[595] = 144'h00faf911ff2f0c51024afa2801e9060d0004;
mem[596] = 144'h0410f43008cd0b8d061c0b9ff8c306290877;
mem[597] = 144'h003beff4001b0953fd30f9c1096701e3fe74;
mem[598] = 144'hf4adf853f71f001ffd090d3505a1fcc404a2;
mem[599] = 144'h02f203dafe6904f5f0b4f6d9ff6ffe2a0406;
mem[600] = 144'h02c80f750556fa5103010027f5abf53ffa45;
mem[601] = 144'h0c75fdd9f171f30107cf09fbfee2f995f746;
mem[602] = 144'h02b90e73f252050a0eb5f60a045afe2ffb12;
mem[603] = 144'h04cc07370e6ffe38fc010c43048cf7ff0d34;
mem[604] = 144'h0d45069400560e1af631f20a0f0e081200fc;
mem[605] = 144'h071bf45ff7c8093b0afafeb208b9f4b8f9b6;
mem[606] = 144'h086104b20b91ef41098f0a2206ca046b0237;
mem[607] = 144'h02eafbbbf48af5d3fb44f546f91b0053fbd1;
mem[608] = 144'h0afbf046f526fd3ef08c080a0259f267f9c6;
mem[609] = 144'hf61df0a9ff98f79cfa3af9cffedc00cbfee2;
mem[610] = 144'hf173fd35f8d1f9a50e14f43508c90212f5a2;
mem[611] = 144'hf4e60635fcc20c98ff320dc6023cf759f4f6;
mem[612] = 144'hfa330cf3fccd000efec7f1f203be0ab1fb49;
mem[613] = 144'hf770f336f4250714f7bbf93702dc0560042b;
mem[614] = 144'hf48b0a50f80df85d066d0b160655f058f8b8;
mem[615] = 144'hf28b00dcfe2701160899f4b107c50a3c086d;
mem[616] = 144'h0744f266f1d907bc020e0e6c019e0414000f;
mem[617] = 144'h0ce504900f3efa4af1f3fe59eff6fffd071e;
mem[618] = 144'hf0e2f64b026b0b4ef15a0e49f56c07b9f8ce;
mem[619] = 144'hf83df9ed05c404b7efedf2a20e38f911ef83;
mem[620] = 144'hfb55098805370cef0c190657f32c00200e2a;
mem[621] = 144'h01ae056109cd030dfbbff7030934f38f0a59;
mem[622] = 144'h03b40660fd620e3f0032f62d0865fa32f2b6;
mem[623] = 144'h09270b07f1870968f42c0ccb0b290992fb85;
mem[624] = 144'h0ba90166fc9af24c0e3c06af08dc05c608a3;
mem[625] = 144'h0e1cfb72fef2f8f105ebf1d70320028df7ac;
mem[626] = 144'h00e6f8180834fc4a0e28f158f485044bf9be;
mem[627] = 144'hf93705bbf7d8fae3f22cf062fc3cf5f9f087;
mem[628] = 144'h0bb707a00c63fb9f04200e65fc8c0308f164;
mem[629] = 144'hf15d0bd3f527fee30457f405f719fdcbf12f;
mem[630] = 144'h08f207e30c1b0e04f2c5ff6a092df10ffb05;
mem[631] = 144'h05bd071a0a64f1380739fcaff1070223f610;
mem[632] = 144'h03320b350402f508f80a04c4fc230c5afdd8;
mem[633] = 144'h05a60e61fb09017afde7f6e5f554f7df06a7;
mem[634] = 144'h0a09fed001d206df01630b860864f44ffc0f;
mem[635] = 144'hf0450712f1a20a5800e507d2f797f280f3e1;
mem[636] = 144'hfc9702c1f980f3d4034b0c9f0239053ff45b;
mem[637] = 144'hfb26fe84fea5f58c019bf83b036a02f80a4d;
mem[638] = 144'h0da60df40da4f761fc7efdaafe3e05e8fb64;
mem[639] = 144'h0c68092507dbf87df0fefe7af2c002d0fd8f;
mem[640] = 144'h0f340c4406a90400f343f00df3fc03b90f8d;
mem[641] = 144'h056cf2b409a10ec9f61c0eca0f2c0dce023a;
mem[642] = 144'hf543f8e6fb9ff6a00d4100f1f0c8f6b601c5;
mem[643] = 144'h034109ba0396f8a80043f896060af4c304a6;
mem[644] = 144'hf44e098103b8068cfee4f1c3f8850f580971;
mem[645] = 144'h07bff322fdc70c4c049af28ff1b6f822f189;
mem[646] = 144'h00b0f4f5ff70fa0c0569f228046ef4b1f5f2;
mem[647] = 144'hfbeaf188fcfdf9e1f76cf2b406aff912ff9c;
mem[648] = 144'hf00e0c4cf614fd5e02b40eb1fa8d0a9b046f;
mem[649] = 144'hfd2b0a990e83f209ff58f31a08dbfa04f689;
mem[650] = 144'h081cfa260800efb6040203fef64f07d2feab;
mem[651] = 144'hfcbc0e2a0e0405d60d250799f2faf08af175;
mem[652] = 144'hfd2d0b9df64503680c03ff400614f92600d8;
mem[653] = 144'hf6540108fdd8f55a0f3cfcd50300fe15fe5b;
mem[654] = 144'hf650f2b903f6051a00b3fbac0ebdfdc6f64f;
mem[655] = 144'hf65a0258f5c40a09f81709130a030d860332;
mem[656] = 144'hf3570e910afefd4af958f7c50d8af0d40af5;
mem[657] = 144'hf765f732f6eaf57a0b8d0a860fbc0f58fccf;
mem[658] = 144'h01f400cef26bfd0af82ff15ef23c0176f382;
mem[659] = 144'h0078fdd9f3600b39f18df930f3c5f438f821;
mem[660] = 144'h0c8cf4ad040df533f58e082df09f0f81070d;
mem[661] = 144'hfdb2fbda06680322f9510a95fd530e380497;
mem[662] = 144'h00e0f23c0105f57307e60243fc3df714f2dc;
mem[663] = 144'h0af5f9dffabcf8c0fc38f918f639fd37fc55;
mem[664] = 144'h0756001b08b502daf4e9049509cd0e280a66;
mem[665] = 144'h0633093f0588fb8f0223ffd70cc9f191071c;
mem[666] = 144'h0996f6caf1e706d2020102e802b80578f360;
mem[667] = 144'hf74303a8ff28fc9af83ff038fbbff309098e;
mem[668] = 144'h0eccf77efa35f73c0af5f77c02b604f4044d;
mem[669] = 144'hf32303d60b51f38ff1acfad10e270399f046;
mem[670] = 144'hf221f92f0dc104a7ff130d33f381016a068c;
mem[671] = 144'hff850dc300fe0a06ef06f87e0f38028df6d7;
mem[672] = 144'hf1af0b0ff91902980a8bf9d504070389f1ea;
mem[673] = 144'hfb29f25006620c87f23bf08df1f6f4330642;
mem[674] = 144'hf702f321fc8ff869059fff98fbf5f8a801ad;
mem[675] = 144'h0f7c01f704ac023df46a07a2f3f2f1530ee7;
mem[676] = 144'h0387f951fb5200760e6afc90067afcd00c6b;
mem[677] = 144'hfbf5f778fc2bf984fd93f588f3010d1e0250;
mem[678] = 144'hfabcf815f393fefff4320becfd3af5bc0e63;
mem[679] = 144'hfb05eff2064f09ae0600fa8ef3810312fa8d;
mem[680] = 144'h07f6f036f247fffcfe5cf5f2f909f0230223;
mem[681] = 144'hfa7f029dfc6100e5f691f7e9f117027f03e2;
mem[682] = 144'h069a057305d0f167f04bf50100bd024e08c3;
mem[683] = 144'hf107fdcbf05bf9d00cf90c98029a0448f44e;
mem[684] = 144'h0542f25f037ff9c2f112faf50e4cf4ff06a5;
mem[685] = 144'hf9c20258fb470a66fdfe0c20f281f1f60003;
mem[686] = 144'hf4f1faa8f1f00cf701b4f4ce0506f2190579;
mem[687] = 144'hfffff3440012f99200340bc4f22b0059ef98;
mem[688] = 144'h0162020d0523f805fecb016efd000563f77b;
mem[689] = 144'h0e1a0791f2dc0b040c98059df0befca6f39a;
mem[690] = 144'hf55afcc60002076bf688fcc90c13f851feb3;
mem[691] = 144'hf241f646fee1f3500ee20bf4f5c300c3fa98;
mem[692] = 144'hf602f20f0438f0650fc9fea1fdf4f603faae;
mem[693] = 144'h0ec7f3990736022ffae105c5f327f1fefe0e;
mem[694] = 144'hfabc01de05aa0bd50a7504cdf61ef868f21c;
mem[695] = 144'h09f6f8920b0dfa7600520f38093f070f0f92;
mem[696] = 144'hf684019c004dfca7fb380adaf6e5fe7dfea5;
mem[697] = 144'h0dbbf499fea6085ef23104c3f57ef264094e;
mem[698] = 144'h042b0be6f187f2b6f0b8f3c005da0b8b018a;
mem[699] = 144'hfb3df3e006e4027f0f0cfd1ff827f41a02b0;
mem[700] = 144'h088e0f350cc5f158fd990baefe59095bfade;
mem[701] = 144'hf3940c21fe3f0ae7f4cf08c90e660174f434;
mem[702] = 144'hf50af8ef075e0d030271090d0840f006f9c5;
mem[703] = 144'h03f8f087febd0ad0fc1e0b6cfd3e0cfdf306;
mem[704] = 144'hfa1af0cdf3510b52f6ae0d3ef1fe0691015c;
mem[705] = 144'h082af03204c80af9039ffd630aa4059609f8;
mem[706] = 144'hf5990346000903bff9d9fd200431fb28f454;
mem[707] = 144'hf996f8d80f7e05d8f01dfe450dee0221f7af;
mem[708] = 144'hf9ff02620766f874f0aa0975fceff1340e34;
mem[709] = 144'hf565f51df95b06d7033e08a6fe49f0d2f02f;
mem[710] = 144'hfa96f3890188f8080ab80d61054aff35f222;
mem[711] = 144'hfb8e083ffac90f82f2450503fa9dfd980652;
mem[712] = 144'hf09bfc6df6d7f7fb0ea0f5d3f0fb05d1072a;
mem[713] = 144'h0ef0f51ef038ff1a03bc0d1a00fe03650598;
mem[714] = 144'hefcef98df55606090e3803c7047f0e100168;
mem[715] = 144'h0df7f108faa6fc8dfad2ff0c070d00af03f3;
mem[716] = 144'h030900d5f784fbf70948f61f05ebf3e302e0;
mem[717] = 144'h0dd6f84dfed7fa98fa690bfbfac7fd3b0efd;
mem[718] = 144'hf5adf29df15a0f2ffecfff47f948f64fff12;
mem[719] = 144'hff8c0686f326f12108bbf550f1e0ef7e01b2;
mem[720] = 144'h095c06bc0fbaf9a203c70603f86906b80303;
mem[721] = 144'h0ebffbbe000dfe8aff6cf811f7690303fe43;
mem[722] = 144'hf54e0082f1dbf51d02b306d400bdfba50706;
mem[723] = 144'h087bf7180419f9d00432faccfd8ff0e8f29b;
mem[724] = 144'hfbcef1a601440644f2c2fd17ffd0f09b0968;
mem[725] = 144'h0cfbfebfffed0dfcfde30951fa3c03180af7;
mem[726] = 144'hf9caf77bfa140d500a9cf60ef5cef60bf983;
mem[727] = 144'h089702670b3cf8cbf79e0247092b0c99fca5;
mem[728] = 144'hf682fec102ebf2bc0e6bfbb5f0dbf466fda4;
mem[729] = 144'hf92dfb2609f507c2f358f5ed05070e590cb5;
mem[730] = 144'hf6050dda031df3d3f897f652f5400af9030b;
mem[731] = 144'hf934f61c0954f8250bbb0297f32d01560891;
mem[732] = 144'hfb58f241f8ecfbbcf360ffb5faebfca6ff51;
mem[733] = 144'hfcc604c60ad3fa56048cfcd2041b0376f27f;
mem[734] = 144'hfbe4fac1f5a6fa7809e1fc19fba3f231f770;
mem[735] = 144'hfa5f05a3f495f3560a1afef4f536fd860372;
mem[736] = 144'hf2480d83f0cafa5c06ca046af3550998085c;
mem[737] = 144'hfe39fd1bf8d30607f00b0af90d1603e603ab;
mem[738] = 144'h0f96fda8059f0bb7fb7d0f2404abf9a204d6;
mem[739] = 144'hefdb060b05690e8006b60e99f86a0c7f0b83;
mem[740] = 144'hf8140770f4cdf5c8087c000dffabf715fc15;
mem[741] = 144'h03620140fe3bf059f0280b990d2e0ccaf3f3;
mem[742] = 144'h0578f4aeff53fd4bfc64f4fe03a9f321f6d6;
mem[743] = 144'h00b20d540802f1daf334f116f09307cb0248;
mem[744] = 144'h0e6803caffd5044ef049f05502aa0e35fc5e;
mem[745] = 144'hefd3095e019cfa8b08ca0691000108fd0a87;
mem[746] = 144'h0e870137efb8efbb01cc0693092f0ab0f834;
mem[747] = 144'h0bb5f43705f6f2f5f5caf414fa9c00a8fffe;
mem[748] = 144'h0138fa57f1cfef97f07dfdc7fcaefb3efdf1;
mem[749] = 144'h0d2a08420a4dffd002380481fb96f7c3ff61;
mem[750] = 144'hff9a0e95f52e0505f6b7fbfc06cc0a4904e8;
mem[751] = 144'h0abdfc860244f78bf608fbd1fb730e03f43b;
mem[752] = 144'hf65dffddff5ffb6108d1f86d04c0f6b908b8;
mem[753] = 144'h031df9f109f8008d0e1601ec0e03030d0f07;
mem[754] = 144'h0d5d0e630f33f611031208dcf71d0ecefd70;
mem[755] = 144'h0e9df51a05d00f3c0e8903980dd9fb520a2d;
mem[756] = 144'h0618f533fd83079e06f80e70f6c50c0a0dc4;
mem[757] = 144'hfb34fa3ffa4cf91d03f70c49f466fbc8f788;
mem[758] = 144'h0b03f1cff4590a70fddff75908e3ffd4076f;
mem[759] = 144'h0843f72cf036042e0adcff2bfba5fac6fa8c;
mem[760] = 144'hf7bb0cea0310f8aa049e0af1077104610e75;
mem[761] = 144'hf590076bf1e008620da1fd38f7c3f038f577;
mem[762] = 144'h09940836f05e03ef07520b71f074f485f978;
mem[763] = 144'h017a0d690ee3efc90092ffa5ff78fe08f321;
mem[764] = 144'hfd660df503cc039ffd990f2c08b606ff0046;
mem[765] = 144'hf07c0da20f88fde2feac00c60761ef670458;
mem[766] = 144'h02b6f6e3f92b0c09f6e3088f01640c190a6d;
mem[767] = 144'h025b08c5ef6b00540176f0a9f33e0294fe9b;
mem[768] = 144'h067f01c1f4b90a070342f039054d0c50fa06;
mem[769] = 144'h0033f4b501e40910f514fc55093ff10af997;
mem[770] = 144'hfec0f415f0d9f53403fff0bf0a9b03400999;
mem[771] = 144'h058401980452fe96f9aff29a04ecfaca0bd4;
mem[772] = 144'h0e3f0dcbf7fa0b590322029e0006fc64f5a1;
mem[773] = 144'h03370587f4630223f155f4effbaaf26cfaa1;
mem[774] = 144'h0da0f8f7f2f40d9ef0820114f3320b5cf4d1;
mem[775] = 144'hf13a04ca0876049e0ded0c940bae0d9e05df;
mem[776] = 144'hef7400b9fb050d12073ffe8e02610a48009e;
mem[777] = 144'hf59c02740c26f5180899079bfff1f9bbfb18;
mem[778] = 144'h0368f6b3f3defb200ad9f58d01e40dd70112;
mem[779] = 144'h0150fb80f3ea0b5c06e207c103950d9f0450;
mem[780] = 144'hf0040d66fa4bf3bd0264f8b1f022f7affd4e;
mem[781] = 144'hfdba004f058bf8c10e4cfd29f51507070930;
mem[782] = 144'h09850e1dfc800e400c17063e08b2081b0f3f;
mem[783] = 144'hf006f526090cfdf00beffcda0a390079ef86;
mem[784] = 144'h0d17f015f3e7f0b3fa910971ff930691f1b4;
mem[785] = 144'hf706007508b10bbf038dff62f895ffacf22a;
mem[786] = 144'h0e69fff201e1f0a904c5f21802e5f93ff3af;
mem[787] = 144'hff7009affd1a0043f047f20b05a906ca04b6;
mem[788] = 144'h0c12fe17049af78c071206170cf4f345f525;
mem[789] = 144'h019dfe38005b0dd3f56ef1ddf387f8ebf493;
mem[790] = 144'hf6e9fd2ef76706ca01610599fff500d7f541;
mem[791] = 144'h022507f0fb10ffd2f594f2d401b4eff80122;
mem[792] = 144'hf9b9f0190123fe020ffafaf8f68707c2ff5d;
mem[793] = 144'h01fe0f33f9520c2705e50795fde1fde400a8;
mem[794] = 144'h06e7f8a2f5c8f8900625f983f2ee0436f11a;
mem[795] = 144'hfd0dff54054c04a7f41901bafefafb2df675;
mem[796] = 144'hf444fbcffd64fdf30702ff410905086cfe67;
mem[797] = 144'hf7caf2700021f77df6a0feebfdc204640105;
mem[798] = 144'hfb6bf6d70c5df13cf2b90626f44f0603f03b;
mem[799] = 144'hfaea0491fac30e0b0066031efeadf1b50c24;
mem[800] = 144'h0ef5feb1fafbf563f7cef9ddf6f30f83050a;
mem[801] = 144'h0622faf4fa5e0a71046604f20443ffc3055d;
mem[802] = 144'h039afbc6f69801300ee7017103d6f51a035f;
mem[803] = 144'h019b01ef017d00a2ff12f0d4f08afeb10a54;
mem[804] = 144'h0147fcccf43cfd820306089e0071f937f2ad;
mem[805] = 144'h022503320cb1fb23f40d00d0f087fe810c45;
mem[806] = 144'h07a70c5f005b0560f7dff3c0f768fedcef5f;
mem[807] = 144'hef99f8070bc004dbfb7bf2dc094bfa7efc6c;
mem[808] = 144'hf52b013af3f205f9eea80ae40aebfe6d0d8b;
mem[809] = 144'h07a2f3b8faf6f8acf50afadaff34fe7f01f4;
mem[810] = 144'h07fafbadf466ff03f794fad1001cfaf804c6;
mem[811] = 144'hf2e1064e00d0f057fece007401e1fe540bb0;
mem[812] = 144'hef28f420f93cf807074305e609de0ab2fb75;
mem[813] = 144'h09d1045cf9ca0511f2e00f500295f0050823;
mem[814] = 144'h0324fe2bf37506f1f130f5940de50e1ef6e6;
mem[815] = 144'hf4260043057a06fdf4d5f294fc5affb904fc;
mem[816] = 144'h07b1f824f0fa00890539f22f0037f1cb0d18;
mem[817] = 144'h04e6ffaa0cb9004b0c3fffc8f958f206f184;
mem[818] = 144'hfce2ff760b84f24a0b5af027f7a4058bf726;
mem[819] = 144'h0bbc0f56f0240510f4680302f6eef3ef0662;
mem[820] = 144'hf093f2e8066b0ce6fce1f4cb08280f9d0c3d;
mem[821] = 144'hf613f9c00d170166f696ff9efa7af5c0faa2;
mem[822] = 144'hfd0f083cf7630115f1aff1820dc6fd08f67e;
mem[823] = 144'hfa8afa34f5b6f1e60852f31c08cc05def1ef;
mem[824] = 144'hfc3c049fff040bfef7cffbbb03c505cafdd6;
mem[825] = 144'h0407fa72fb12ff25f584f6c7f3df051ff131;
mem[826] = 144'hfe10f9120496093e02a6fc1ff2bbf78bf5df;
mem[827] = 144'hf2090cb00e8af95a0884fbd7098efd59f018;
mem[828] = 144'hf86f0145f05dfa0bf941f1f2085dff5d0b29;
mem[829] = 144'hfa440e89fc36010e0c6a07b10083013df6a7;
mem[830] = 144'h0d6ffd0df20bfb93f663f11a0f4df2f4f2a5;
mem[831] = 144'hf81002f0fc400c3b025900a2f5c1fe0ef960;
mem[832] = 144'hf4a10b0efd6ff133ff5103850f67f257fe43;
mem[833] = 144'hf81601b6059df2ec08bdfddaf201091a049e;
mem[834] = 144'h0a46fec4014cf08bf183fcfa075800f20e01;
mem[835] = 144'h09f0fd3b0c67f505fb5f03faf8590b970607;
mem[836] = 144'hf20df023fcbff2d1fafd01520e8903c8fc99;
mem[837] = 144'hf699f1fc0f0a08f1fdfe0c790edd0c32f004;
mem[838] = 144'hf1b00d2f024104ce0ce20179fb4a08bdfb4f;
mem[839] = 144'h006ef474fa780d5a0aeef0b70c110ca00d0b;
mem[840] = 144'h0b15f4b1f910f215f0d4fa240082fd4502e1;
mem[841] = 144'hfaea0b4df27c003cfda5f872022b0b3400db;
mem[842] = 144'hf582f2f80bd20dfef60b051802e6f6b7feef;
mem[843] = 144'h025505ce08510352f2c70ccb02eaef69f5c1;
mem[844] = 144'hf01208b9f818fa68fe7b0362f85c0d9403c1;
mem[845] = 144'hf4cf0ec5f9d70ac2f8950245f238044b032c;
mem[846] = 144'hf892f567fd98faa706da0f9a0f570b03f850;
mem[847] = 144'hf670ffb2f04904d100ccf3c6081d0f48f690;
mem[848] = 144'hf4edf1ea0208fa690181f51c0936efc10044;
mem[849] = 144'h0b650269028d055d07c9fc420549f29108f4;
mem[850] = 144'h0796f04d009af0b8fd61f54cf51df445ef4b;
mem[851] = 144'hf17f09490e67fbd4fe850c13fa6a056b0387;
mem[852] = 144'hf8b1faa207980c6cfa78f241f7e6f1900536;
mem[853] = 144'h0ea7083fff5508460ec10a6af85cf260fec4;
mem[854] = 144'hfc3d097dfcbbfbb2fd980605f55c0cf807c9;
mem[855] = 144'h093908710ce709a8ff530daa00a40938fd43;
mem[856] = 144'hf8c20e11fcf807450901039d0193ff700c94;
mem[857] = 144'h04ab06eff6cbf28306120439f9e30d8f09c2;
mem[858] = 144'h003df2e100e90fd40dcc04020beef678f863;
mem[859] = 144'hfc4c0899f983f6abfe6bf059012ffd960878;
mem[860] = 144'hf7b1fc370496073a02040fdd0a8df7960888;
mem[861] = 144'h0edd0e09f47bf761017cf489fadff447f93c;
mem[862] = 144'h07e604a70d54f3990d62eff10ec70bbfefc8;
mem[863] = 144'hffa9febc08bff2280235f2ee099107e00be7;
mem[864] = 144'h0ce40de7f733fa970e04074e04530c340caf;
mem[865] = 144'hf7a70c4cfd950b15fd71f8bd07b8fa12fb8f;
mem[866] = 144'hfdc3f799f7c5f7d50a47f29409a60bda0d19;
mem[867] = 144'h0cfafafcf63f099ff13d099dfcc107070d4b;
mem[868] = 144'hf8a9f5db0d72f8c1f62a0434fe76fe9bf4bc;
mem[869] = 144'hf6ae00ad070f0a2701850d4ef469fd77f816;
mem[870] = 144'h0483f5270d73fc06f6f201a70b6f077d0fac;
mem[871] = 144'h0647ff90088203e1f30e0f25025e0c3df12d;
mem[872] = 144'h0690095100faf3d004d204ab0bc7f0280d69;
mem[873] = 144'h08a6f88ff6ee08170a7503a0f11df95b01cd;
mem[874] = 144'hf837f9b9013b0843f57df9e6f176fdfa05ba;
mem[875] = 144'hff19fb82f929f543075efb810028fbc00e47;
mem[876] = 144'hfb08f408fca7f08bfb9107710554031c016f;
mem[877] = 144'hffc5fd5bf622f593fdca04d105d001a00a78;
mem[878] = 144'hfe2e01a7f6ea065cfd1c00290eeb019e0eae;
mem[879] = 144'h0ed50221febe0e9e06b5085400a6f4a3f016;
mem[880] = 144'h05620d77034b08bf079aeff904a1f1d9f0e8;
mem[881] = 144'hf8ecfeedf74cf057fe68f1a6077cf21df175;
mem[882] = 144'h018efc17faad044af63ff6e60035025cff2b;
mem[883] = 144'h01fd01830ab60207fc140e19fe800bf705c9;
mem[884] = 144'hfc8ff37ff3880e60fdea094ef7f1f70afe6a;
mem[885] = 144'hf655fba5091f0d10f2d1076b0a16f390fe03;
mem[886] = 144'hf0b2fbf30ac40d1cfeb90bf3fe960b020687;
mem[887] = 144'h07a70443fe8404630191f8f90690f16df422;
mem[888] = 144'h06d1fb84f137f172f37700b506370337f7b0;
mem[889] = 144'h0893f74afd500d7cfcd10f46fe9d0a0bfa6f;
mem[890] = 144'h03a2f601f7e2f794fd95f340f0cbfd190cee;
mem[891] = 144'hf85908bcf003f047f5d0f16ef46a035c0071;
mem[892] = 144'hefb7f8b2fee708d706f30772028ef63ff329;
mem[893] = 144'hf249f16ef0e4f866fcb307230e6501dcf7bd;
mem[894] = 144'hfb09ef82040600a9089df4860e4cfb890c39;
mem[895] = 144'hf244f3e409b5096ffa55f555f204f5a205cb;
mem[896] = 144'h0ce7048cffc6fb24067afc3af3ebfd020910;
mem[897] = 144'hf8c0efebf2ff0f790523003d05e702330948;
mem[898] = 144'h0387f105013c00c7f961f6b70411f2c50338;
mem[899] = 144'h0d6cf5820475043e09b50106ff4efc4deffd;
mem[900] = 144'hffcf0fda0efa0af5f982f927025a06cff1ca;
mem[901] = 144'hf1d2f433f235fe0e0861f05f0baa0a0e042c;
mem[902] = 144'h0185fea50f1701ebf3ce062dff0cfb7d00c7;
mem[903] = 144'hf7310786034200d2f2cdfc2e0bda077c0e08;
mem[904] = 144'hf24efd03fb740cad002c01ea0070f83bff9e;
mem[905] = 144'h0263f7c4095a0daf04af095bf9a5f859f456;
mem[906] = 144'h02e80569fc6d0e6007def3830328fba4fa73;
mem[907] = 144'hfd940008fbae0ba403d1f24f0f80ffaf0a00;
mem[908] = 144'hf4d5041d073d090eefc50e870aa60c96f3f3;
mem[909] = 144'hfd8d02cf0f6100d1f1860a1bf8d9012bf597;
mem[910] = 144'h089afb86f02f00ee07270b36006cfda3053c;
mem[911] = 144'hf923f184065c0d560a73f1420a6e02100262;
mem[912] = 144'hf9ac07cb0b7ff995fdba0674f2e3014704bc;
mem[913] = 144'hf0060b4705e901a4ffebf0cffbb707ff03e8;
mem[914] = 144'h0791ff540aeaff990060f728047d0465056c;
mem[915] = 144'hf7430876f96f0602fbc1f7660880f74406fe;
mem[916] = 144'hf29902cef1e0f7f50bc3fb3301a209ccfcfd;
mem[917] = 144'hf977f875f17d06b5f69408ae0409f43cfcc8;
mem[918] = 144'hf28c015f0bd0f584f26107b30053f08305da;
mem[919] = 144'hf4eb01d1fb2d0360f2f80203f222fbf0fe45;
mem[920] = 144'h007e0582fd2200eb0e09f7ec0d2cf4f005bb;
mem[921] = 144'h0761ef5ef8f5f10f0576f0b8041dfb2201ec;
mem[922] = 144'hf4370cbef98ef2290609076dfa32f82e0ee7;
mem[923] = 144'h092df3510f42f2150afcf8d8fc38f0d8faf3;
mem[924] = 144'h08b5f7a8000efa7b005a0ad3f6c50ba000f9;
mem[925] = 144'h06b5f554ef36f89801e1f2e1fae50371fe86;
mem[926] = 144'hf8d1f120016e0ac70f84f3f1fc53f539fbbc;
mem[927] = 144'hf85103d0078ffcb1f64308850d080c7af9d7;
mem[928] = 144'h059d00d907a6f42ff5c5f74d0296f4e9002c;
mem[929] = 144'hfdfe0f64004bff5bfc4cfe7300f008470919;
mem[930] = 144'hf774fea603a20bb8fc84fe760a20f5b90a19;
mem[931] = 144'hf6b9f79e01eaf0d6f7020ea0fda8eff80473;
mem[932] = 144'hf98cf6d1fb650112ff5bf7ee0214fe650c56;
mem[933] = 144'hf2eb0de90b3f0f46f80d06e8f4a9fe630c43;
mem[934] = 144'hfc8cf5c3fe2b015e090802660e1d02f6f8de;
mem[935] = 144'hf656f774fb0302ccf9d903d909c0ef87fe9e;
mem[936] = 144'hf572060204a0f99302bf08d60654f1aa04e1;
mem[937] = 144'hf7e60521f06000f3093ff8d8f8b4ef53024a;
mem[938] = 144'hf94c0485f57505c50433f60af24505850975;
mem[939] = 144'h07180a900743f9c5fac9f43401e7011c0d1c;
mem[940] = 144'hf53af0970a57f0dd04d1ee74f138f0d0f5b2;
mem[941] = 144'h0155efabefd7fcb80657f15af22ff765096c;
mem[942] = 144'h01080863049f0275f8ecf726f430f59d02dd;
mem[943] = 144'h0aa6fcacf6700a88f11bfc88049afcfc0233;
mem[944] = 144'h0b5b08fcf4cd03e70cd2ff39f84b0d1b0af7;
mem[945] = 144'hf893f0eafac8073f0e8e0fb30ecef6c70bde;
mem[946] = 144'hf89b0834ee4c0a4c0b1204e1ff4c002df3bf;
mem[947] = 144'h0354f63602ca0f04ff38fef80d5bf00206ee;
mem[948] = 144'h0eecf28ff1e6f113fbe006c2fa39ff05083f;
mem[949] = 144'h02f9087cff7ffd4909cdf372f091ff6ef53a;
mem[950] = 144'hf0ac089dfc4a09820227089bf8230f8ef8c3;
mem[951] = 144'hf0de01dbf3210a34fa87f6b2f3aff7500242;
mem[952] = 144'hf6b10b4f0248fac90ec30c4903980e6c036d;
mem[953] = 144'hf395fb53eff9fabaf5de0445f709fe3f0d4e;
mem[954] = 144'h0eaefe8ef3da01330972017ef023f191f394;
mem[955] = 144'hf268ee6a08b6fbb2057dfa1df31cfe780374;
mem[956] = 144'hf5adfb4ef1d0fd9cfe230b020c520c2b063c;
mem[957] = 144'h0b2c0a9bf0e7f42df480feb6030a0dcef11b;
mem[958] = 144'hf96a0ec1ef6705c4fc39094105d20c1e050e;
mem[959] = 144'hf54d05e0063df27208eb0252f1f6f350f298;
mem[960] = 144'h07f7fbf1f506f88e076bf42e06890914f0d4;
mem[961] = 144'hfdfafd8f0bff0ff3f4010ee703cc03520e5f;
mem[962] = 144'h0e06f1e60727fd07045df7f90871fbeef431;
mem[963] = 144'hf8c40b53f21d0cc2014f018df138f9a708d1;
mem[964] = 144'h04c503d5079005860f6dfa4b075904280d38;
mem[965] = 144'hfa41f62afaa7fddc0c90fa2bfc49f4b1048f;
mem[966] = 144'h04aa022af7b7ff0d08310db0f093049d079f;
mem[967] = 144'h08a10387f4740cff044502b10f190cd3f8b1;
mem[968] = 144'h0f37fd07f600f5f30caa0c12fe680127f56d;
mem[969] = 144'hf8fcf431fec30c790658ff7cfe44f9d3f3e7;
mem[970] = 144'h008d0c2e01ce09e4f40af745f7580e9cffd2;
mem[971] = 144'hfbb1efd20421f00df45907e2f415f3fe01db;
mem[972] = 144'h02fd01d203f70aaaf47e0017fa18f5b5f88f;
mem[973] = 144'h04740039f48dfb1e0bf20fc70228ffb4f4e8;
mem[974] = 144'h0f240499078607f5fcda0aeefcfdf2b600c1;
mem[975] = 144'h030dfff409be09830d6d08f80ca9f7e406c7;
mem[976] = 144'h0383fae200bffa6ff6ebf61a03d70b0908b4;
mem[977] = 144'h0f6af6010556f96003170b050978faeafdfd;
mem[978] = 144'hf8b0f46befcb013805a30d3af682f8c2fb40;
mem[979] = 144'hfdb4fa620c8101fcf3e00c1e051e074f09d9;
mem[980] = 144'h0bd40460f2dcfbf4f98d09240e65f67308e0;
mem[981] = 144'h0568ffd102c0f63002820da003a0f2b0f294;
mem[982] = 144'hf95dfe56f1db07120e42f03700120aeb00b8;
mem[983] = 144'hf2ccfea2f062fdf9f907f7d709d8f9acfed4;
mem[984] = 144'hf8b70c780245fc2009cb06ddfe53f72f0e95;
mem[985] = 144'h0008fcedffd0f1f305c201c60679f8bf089f;
mem[986] = 144'h020df2f0fb5eff5408270862fa53fe61f2a5;
mem[987] = 144'h05400342f33afd8cfa8d0579fa280025fe15;
mem[988] = 144'hf8ddfa250b020917fbd8efe408fc01b8f993;
mem[989] = 144'h0d6c0d9dfaaff274f3c20a370f050230061c;
mem[990] = 144'h03610e2804620ea0f03af0aaf058f259f5c7;
mem[991] = 144'h04060b460379fd6afcbff035f70ef928f15b;
mem[992] = 144'h02a40714fe33f45d0d4afd6f0fd6066005cb;
mem[993] = 144'hf128ff19f043ff1d0e60f05df515fc58fb91;
mem[994] = 144'h0dc0078b09500e230420fa38092b09f003cb;
mem[995] = 144'h0a4ef15ef25bfad40cc1010bffe8fb13ff59;
mem[996] = 144'hfc1d013b007c0c210abff3fa0727f63e0c0c;
mem[997] = 144'hff2ef46dfb6cf7aff7aa071eef76fbd2074f;
mem[998] = 144'h07db03670344043609dfff8ff029f0c80610;
mem[999] = 144'h0042fe89fbf5fe03f9b8f3560b080c0d06a7;
mem[1000] = 144'hfae0f1e909fbef540534f257f7c806400ec0;
mem[1001] = 144'hf6d00379033c0c0afd6dffa3fb990a20f0f0;
mem[1002] = 144'h074302150b95f972f243fc180601fcc80d5c;
mem[1003] = 144'h08100908f6a60aaf0ccc0c52fa30ff53f022;
mem[1004] = 144'h06b6f2c4ffe3f5c8ff17f5e1065fff05fd0b;
mem[1005] = 144'h0ecdff8bfb15f874f5f8f8e50e92075cf5f0;
mem[1006] = 144'h0badeee6098ef193f59ff8600874f81ff1bf;
mem[1007] = 144'h082e08ecf5a7f0b4efcb06a8f5d6ff9d0e3d;
mem[1008] = 144'hf3daf8600647fe6df218f3d4f7110e7ef1bd;
mem[1009] = 144'h0b290492fe0cff7e04abf88afdf405cbfede;
mem[1010] = 144'h0aebf6d2fc440b0dfab306acfcca0d5bf0a8;
mem[1011] = 144'hfc84ff1a08cdfcb8f4d4fcde01aefc480645;
mem[1012] = 144'h06f601930e51f5be096cfd8a089cf54bf4f1;
mem[1013] = 144'hfeaff4390b35f60507cef22beffb06bceffd;
mem[1014] = 144'h0f2cf596f68207c5f70702490a3dffdb0449;
mem[1015] = 144'h0580055a08b90a040d1008600bccf8020b2c;
mem[1016] = 144'h05710e09008104eb0e9bf44bfbf70d480ccd;
mem[1017] = 144'h0e4e0b77f7350dfc05a5010b04750d27f412;
mem[1018] = 144'hf58d074f076209b5f0ea010407ea0b2df22d;
mem[1019] = 144'h0947f9620c01fdca07b7f7f00557f1fff462;
mem[1020] = 144'h0415f46e04d6025bff14ffbf09cafb3f0266;
mem[1021] = 144'hf924f3a7f999fd3eff0c00a907c6fb63f519;
mem[1022] = 144'hf1c006aa05ff0a15f0b5f979fc8f009d049f;
mem[1023] = 144'hf03b03affeb4016ef6b10a36f309f168f724;
mem[1024] = 144'h02470f83013008f9030f0d3dfc7dfcd30e86;
mem[1025] = 144'hf0160d9dfaef0919ff54f396fcfe04d0f1a9;
mem[1026] = 144'hf06a0a9efcb80918f630f69501ca0649fd3b;
mem[1027] = 144'h060506bdf913fd5dfc39007b0a34fddc0f21;
mem[1028] = 144'hf15af0f5efd80c59071bf0000edf0de80b5b;
mem[1029] = 144'h0d01017f055ff3810760f81eeffb0f58f290;
mem[1030] = 144'hfdb9fb3902acf4790809f4550345084f080b;
mem[1031] = 144'hfdbc098efd6ff2d2fbe607bcf940f81f06ef;
mem[1032] = 144'hf52e0d12f26f0e20f032f5fcfbdbff5b098d;
mem[1033] = 144'h0802f62306e5088c073405e6f0d1fbd9fd0d;
mem[1034] = 144'h048902020bf80076057cf4b5f6d003cff0f4;
mem[1035] = 144'h09bb0ecb0b97fad4fa0601eefa43089ff9be;
mem[1036] = 144'h0a0e048afcf10623f853fb2efcbd041af825;
mem[1037] = 144'h0856f513fc950ed803aff7a40e1dfd71f443;
mem[1038] = 144'hf16ff6d00adf01f60b1a0c67faad0e62fe51;
mem[1039] = 144'hf1a102de039cf23afc4a0c700c77fe3e003e;
mem[1040] = 144'h0d38fd66f369f5fcfeaffc48001dffecf071;
mem[1041] = 144'h03f90df30681ff83050e08f6f7a5fccaf4da;
mem[1042] = 144'hefdf01c90dd8087703b007eafa66018c0db7;
mem[1043] = 144'hf43e0e210dfe013ffae8032d053ff540f812;
mem[1044] = 144'h026efcec01d9081cf34107bf0438f40802a1;
mem[1045] = 144'h0ef4f00e01a40867f183023ef0800d57f88d;
mem[1046] = 144'hfcc8fc06004c01b5fc5c0ac9f703014d01ca;
mem[1047] = 144'h060fff790d8aff8305f3f66cfa740502f934;
mem[1048] = 144'hf23afffe05faf83f0a58f9b7f78efdd90864;
mem[1049] = 144'h0e540edaf1daff66f70af4d9feba04ef0470;
mem[1050] = 144'h05c8f274002afa6f09ea0894f1acf53d0e51;
mem[1051] = 144'hfe16fd61063d0303fc750658019b030df908;
mem[1052] = 144'h0bcc0b3f05cdfe6c0489057a08b50733f510;
mem[1053] = 144'h01faf67cfd1809a10eabfad0f90100690c93;
mem[1054] = 144'h04b7f8f808a70481f4b5fa2afe85f4da0a86;
mem[1055] = 144'hf7fa0bb4f9580986f5a6f04702a200110a85;
mem[1056] = 144'h057cfd58f75cf38406b10bff0d7bfc38fee8;
mem[1057] = 144'h076bf30804f405fffff8fd57050e027808ff;
mem[1058] = 144'h042103ae048b0a80fc62f03c09d905b0f3eb;
mem[1059] = 144'hf0740f8807410d0f03060a3a0314f1c90d51;
mem[1060] = 144'h0a8c0921f9b70541059e04ecfa23ffd1fcec;
mem[1061] = 144'hfbabf3b4fabd0f6c000f00f6fb45063b069e;
mem[1062] = 144'hff44ff37082a0cbc003305b3fc5f0b900d8d;
mem[1063] = 144'h0cf8f568f6d70163f34e06d8f50608e4f501;
mem[1064] = 144'h07adf0f40924f8c1009ef0dcf782f36b0d43;
mem[1065] = 144'hf3a1f9d3f8da00bf01eafe8d0d84f0d5efab;
mem[1066] = 144'h02c90bcd01670084060e0c770259f1ae04ad;
mem[1067] = 144'h0da8fbc20229fbf9faebfe3cf2defe69f3da;
mem[1068] = 144'h0a3d09cefb8b04cef089efb2f73e0aa102f8;
mem[1069] = 144'hf5b1f337f3d107bd0ce2f384fcdc08c0f0a3;
mem[1070] = 144'hf8c6f90b0aa5f539002af3f4f9b6fc97083c;
mem[1071] = 144'hffcdf3b70090041301cffa24ff6606580b0d;
mem[1072] = 144'h06db0f3ef7830f350c41fffb05ebf8ac0ddb;
mem[1073] = 144'h04c6f34ff28ff5fef9fe0619f4e5f78cf56f;
mem[1074] = 144'hfc1ff03cf3a5f21f0f55059c0c030a34f7c1;
mem[1075] = 144'h0d53f5e909c4ff64f83f05ca0d85080e0d0e;
mem[1076] = 144'hf56405d5faa401560a690ab2f1a7fe2d0631;
mem[1077] = 144'h08b9063bf987ff8dfe01f07f00de04ebf0bd;
mem[1078] = 144'h0ad6f962f3ce0e64fac7fda8f13ffdc1fe57;
mem[1079] = 144'hf8720bc60a70fad3f6c90d90075af0b4fe86;
mem[1080] = 144'h047907600dc40a9af7330280f00606b10b08;
mem[1081] = 144'hf4d7efc3f122f211fe7ff923fab7f9c30ef3;
mem[1082] = 144'h070ef3acfa3bf7590786020afe0e08b60a81;
mem[1083] = 144'hfa34ffe5f18ff33ef67201490a2702e60bb1;
mem[1084] = 144'h04e8fd81fdcdf528fe4a0a4d011bfe430067;
mem[1085] = 144'hfe400c24ffa2f1dafa29ff680308f0aff635;
mem[1086] = 144'h0f000bb6009f0d79f6a6014efb4df496efad;
mem[1087] = 144'hf5db02a2f6b3f35ef70804d001a60f2bf6f2;
mem[1088] = 144'h06f4060103600d0a01c6fdfa0ab0f41a0f8c;
mem[1089] = 144'h0f3c049af538f37d02fff7080c740593ffb2;
mem[1090] = 144'hfbd5043a04c2058af30afb81f77904ac0151;
mem[1091] = 144'h0bd70434f345f56406df04ff0245f1810a0d;
mem[1092] = 144'hf997000212abfb410aaf0b82ff13ff39fd1f;
mem[1093] = 144'h00650787fa8ff2c1f08cf6c304b304670e5a;
mem[1094] = 144'hffb2f2df0e11008cf0460c25f0fa028b04ad;
mem[1095] = 144'hf1a006cc0be3f5c4f32af1b8fa04fbf4fc67;
mem[1096] = 144'h0bb7026807f9ffc9f7eef3890d2702fefe4d;
mem[1097] = 144'h0cf5f45ef794fc0ff6eff4dffae403b6fbf7;
mem[1098] = 144'h01c90a39ff13078204aafdc9ff89096f0e47;
mem[1099] = 144'h05b4fb38ff5bfde5f7b6fbd5f7c8f985f91d;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule