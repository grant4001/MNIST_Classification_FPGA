`timescale 1ns/1ns

module wt_mem5 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'hf735f30af566fb7206a5f5b5030d04e5f050;
mem[1] = 144'hfea20768f0130bb20332028afecbf50b0ecf;
mem[2] = 144'hf27cff5bf91b0e2e0a58fc79f0120c200ed3;
mem[3] = 144'hf66dfe4a0ad4f5730db8fe220650f839008a;
mem[4] = 144'h034ef3070396f8c60b48f43603960820f059;
mem[5] = 144'h0b74fbd3fee3006afe6af2c80322f8baff19;
mem[6] = 144'h032e0b8efac4ee7906920691007df442f9ea;
mem[7] = 144'h0c8903def70df8210a15f737f0fcf64bf8ea;
mem[8] = 144'h0b560c96f6d5fd09f0b0f71df1b2086cfbd6;
mem[9] = 144'h0d700746f07401a10b3ef7dc041afb1efd0d;
mem[10] = 144'h0c6d0aa0f8affeb3f73d0015f32a0c55fb91;
mem[11] = 144'hff5702de03a009150b2d0ae205cbf6ed03a8;
mem[12] = 144'h00ab01e704860b58fdf4005f0810f9c3f9f7;
mem[13] = 144'h026d04b7fe13f6f3043f06b80bc8f070fbd1;
mem[14] = 144'h0a28f3f10cd6051efa700362046b05f7f9d2;
mem[15] = 144'heeef0a7f04020439fcbafc4800040d1cefba;
mem[16] = 144'hef9b0cf706970937f36d04ebfc6fff02f8a4;
mem[17] = 144'h0743026dfd88f4e8f75fffd8f80a0883f56b;
mem[18] = 144'hf76af214eef2fdf3039ef5f4fa3ffe4706f9;
mem[19] = 144'h0268f561f579ff5a069a0e1304170142f0aa;
mem[20] = 144'hfd3bfd18f048ff50f2edfd790497015b066c;
mem[21] = 144'h0532f212061d057c006ef79107f5ff3cf7d4;
mem[22] = 144'h02cbfc4c01ef06d7fb0404f6fb1f016efa13;
mem[23] = 144'hfc5bf132fb3805b20907016d0a4dfafeff3a;
mem[24] = 144'h04b602f2f95c0ce0039f0cfc0d3305620bdf;
mem[25] = 144'hf05f058d08ccf4620729fa7cf6ef0a310466;
mem[26] = 144'hf3ae07b9fe500aebf4cb061efb0a01c4fc86;
mem[27] = 144'hf3610d8d081bfffcef3efc5303acfbc40083;
mem[28] = 144'h0dd20648f0b3ffcf0da10b7d0287feeb0012;
mem[29] = 144'hf508fa88ffd6ff9ffc2a084805c0fc090e34;
mem[30] = 144'hef75f0d6f7c2f81a028a0ca504ee0b28f847;
mem[31] = 144'h0d31f206f3d40cce0c68fbeb0d0ffd690bdb;
mem[32] = 144'h0ba5021bff85f540fa12fcf40670f45105ba;
mem[33] = 144'hf5f9f160074bf0990591f2a00ba7064df91d;
mem[34] = 144'h0a4e02b70e3003410d7808110e0809e20c17;
mem[35] = 144'hf6c1f47ff6afff9bfceef748f52bf4e80573;
mem[36] = 144'h0705087bfa60f839fd2ff9a5ee6b09eb0834;
mem[37] = 144'h0e74f8a6fcab0ef90b38f37f050cf41e0ab9;
mem[38] = 144'h01a00d22f7d1efdcf910fe37f66605b30195;
mem[39] = 144'hefb002c20d4b0a85f7a908aefd8f0c88fe65;
mem[40] = 144'h096bf6b4f037fb41044703740836efc1f80b;
mem[41] = 144'h0f57fde50286ff90f7e9fa520c7dfa280380;
mem[42] = 144'hf1450200f27afce30f2e0572ff4cfba9f7d9;
mem[43] = 144'hf2810d2dfa9bf791f83c07450d40fdf0fbc1;
mem[44] = 144'hfd54f66df557f288f1e8f14bff09f0110d80;
mem[45] = 144'h07beef98fa4d05c20d81029808c1081102b0;
mem[46] = 144'hef900b99fb800e35fc5a0929fa6cfd01ff2e;
mem[47] = 144'h0c7b061b05f206bef73dfdd703a70d9e0efe;
mem[48] = 144'hf483f24bf0f1fb41f24e0b72049d02d8f373;
mem[49] = 144'h09faf40bf5bfef36ffbcfd650e3cf434eeeb;
mem[50] = 144'h011afe2a09ddf46eff73f6500bbaf86207f0;
mem[51] = 144'hf8ee031ef774f104f604ff810020080e0e05;
mem[52] = 144'h0d35f78801b10398010ffda0ff5a0c26002f;
mem[53] = 144'hfc70f61cf658ee890a67f858f0090a22f043;
mem[54] = 144'hfcbef9acfd790e7f0f41f421f38006440901;
mem[55] = 144'hfa4207260031f397f5c504500738ff2c0876;
mem[56] = 144'h0b29efd502d1f54bf9cef993ef2afc2bef85;
mem[57] = 144'h024bef96fa66f07dfe82f93205faf385fa7f;
mem[58] = 144'h022ffe39f7200cedf3e9f6a7011dfc1b0f02;
mem[59] = 144'h052a015df7cb0f5c0c9cff0106fff37bfc27;
mem[60] = 144'h07a6f45dfd1307a90b0dfb450d86001f0889;
mem[61] = 144'hff46f46cfc4c023e073af6aaf0adfe5afc39;
mem[62] = 144'h0b03f48cfaff02c0fb15ff190de0016aef66;
mem[63] = 144'hf7ba0573010bf4e301ad06da0cbd099d04d9;
mem[64] = 144'hfe0df9a3021f012ffab804bb022ef7ad052d;
mem[65] = 144'h084ff889f47af314f9fcf211f90508160803;
mem[66] = 144'h09e504020032f66e002a0ba9f01709a0fc85;
mem[67] = 144'hfe42fc7a0ae2f2540420fcacf20203ea0c44;
mem[68] = 144'h08fb0011ff17f0c5f969084c0bf300a30911;
mem[69] = 144'h00b5f80cfcea012c0e040181f127093f056d;
mem[70] = 144'hf8e50d11f850f4460d5a0b5dfc69f38d0b47;
mem[71] = 144'h0cfef5c4fefaf64df667f4d1f562fa0a02bd;
mem[72] = 144'hfa370cd40cdffb12fe05fbcff85e0174f280;
mem[73] = 144'hfa3d08fff8b1fa13ef3e0ce50b6af27c0a8b;
mem[74] = 144'h0cec00f8f809077f038ffc830187fd44fa99;
mem[75] = 144'hf35d039705f5079703130a2a0b51f544f15a;
mem[76] = 144'heed9f5fcfae1f2150ba1ff49f1970134f699;
mem[77] = 144'hf79b02f10aa10d980b7aefc90ed30141fd3e;
mem[78] = 144'h0a730a38f47bf407039af16ef14af7920243;
mem[79] = 144'h06dbfd250e3d0a660957f6b8f982006af4cd;
mem[80] = 144'hf13a0e32fde401a60c5df34af9eff163f856;
mem[81] = 144'h083703fff379f2c7f4320bb60bbd0d5ef6d7;
mem[82] = 144'h00610199fdb4f31106e001c0f2750a5c03f5;
mem[83] = 144'hf0b5faf10a360a1cf4f001f3029ff5fafaac;
mem[84] = 144'h0e27fecef43ef3acf1990a63fc9efb65f706;
mem[85] = 144'h074cf303f0b70e6cf7d8f841075506530369;
mem[86] = 144'h03baf24cf33205690864f62f0ba503de0e23;
mem[87] = 144'h04dffb5b0f22ffb2079ef4530e2cf8cb02ce;
mem[88] = 144'hfdbcf131fd550ef9f076ff2d0e5ef68100b0;
mem[89] = 144'h0e1e08ccff730ab003cfeff5083cf0fc0399;
mem[90] = 144'h05280095f02703b8f06fff640ba70461f545;
mem[91] = 144'h06990278075608eaf8ecf618f1c20d96fe28;
mem[92] = 144'hf47d04d7f21903cf0c35f56d0ed1fd640edb;
mem[93] = 144'h04f4fcbdf8bc0f1ef919091ff3a4fc7ffc58;
mem[94] = 144'hff54090dfe1e042207510bb0fca0f64bf18a;
mem[95] = 144'hfea1072b0652fd87039302ad0651054209b2;
mem[96] = 144'h0e6f03e6fe6e0b58f5d2f6ddf390f18ef953;
mem[97] = 144'hf856fd8d091bfab1f71af9060423fcfcf5af;
mem[98] = 144'hf95ff679043bf4ac061503a807f8014c01df;
mem[99] = 144'hf6b602ea05e3f3310787f0e1f907fcdaf064;
mem[100] = 144'hfe2a0ade0c260279f308f012fabbf13bfc61;
mem[101] = 144'h0044f840fc6cf8f809650787fed9f081f5ad;
mem[102] = 144'h0a6cfd410d8bfe2af7c40f0102f50085fd06;
mem[103] = 144'h09ff00fffcb60202fe4402e2f4fcf01afa05;
mem[104] = 144'h0d220c88fa5905f006e109cdf2310835fd82;
mem[105] = 144'hf10df4d00a13fb4e0d200c4d0250fd8d01b5;
mem[106] = 144'h01ac0181f56205550becfdaefb500318ff3a;
mem[107] = 144'hf4c40e1e0b7409c6fd2907d2ffd1f717f2d9;
mem[108] = 144'hfdd8f173fb98041801a7fd95f6d0f366f327;
mem[109] = 144'h0a58fdbff533fb1bf37df752fb94fd0df043;
mem[110] = 144'hfc7c092ff119fec508bdf2f2fdbcf08ffac0;
mem[111] = 144'hf07afbb0f425ff50063d0b3ef596061d0bd3;
mem[112] = 144'h062df8d2fb85f12b066a0efaf0d205bff840;
mem[113] = 144'hf852f7760a6407410f75f488f604f677fdef;
mem[114] = 144'h0893fa3e084801f30485ff9a075001280383;
mem[115] = 144'hf27df96b086bf7d004e90ea10c77fbdcfe04;
mem[116] = 144'h0d7e05eaf76bf290f5dbfcb006c5ff0c0731;
mem[117] = 144'hf4e70afb068a0b1df0e40568f0e6fce0f32b;
mem[118] = 144'hf958efe7fe510b060573f2250a4cf94809cb;
mem[119] = 144'hfab604a90885f95ef153fee20d5cfffef038;
mem[120] = 144'hf5b4f35d0c78efea020906c80df2f9a503eb;
mem[121] = 144'h0ab50b15f8b7f433f368085507e5018400bc;
mem[122] = 144'h0140f6b4018df14df97ef53ff58bf14f07ce;
mem[123] = 144'hf3e3f3fef3540688079e013f0e850792f6a4;
mem[124] = 144'h0e1b0b03f0d8011bf478f4490f21ff94f804;
mem[125] = 144'hf5c8f9e0080f0ce90dd2f52b0df2f97ff154;
mem[126] = 144'h05b60cf2fa6ff416fbdd08faf8b60b4c06fa;
mem[127] = 144'h0d3008460ccf0dabf229034d07e4f7dc03a6;
mem[128] = 144'heff0f44f0350f568fbac094c0e04f03a01e1;
mem[129] = 144'h0454fe06fae907a8fdcdfce904af06b90292;
mem[130] = 144'hf24008eef9c70647fe82f735fe3c08390b70;
mem[131] = 144'h09b9f0bb05f3f54f02fbfbdaf3b60b100c15;
mem[132] = 144'hfdbef466fbbefbbdfd2504c4fca6fd2df6c0;
mem[133] = 144'h098f0950f59df3bf0ec3f7910a34f63dfb37;
mem[134] = 144'h0c9d052ef9970a8500d90ddf0a76f23a077a;
mem[135] = 144'h01bd0653fbb00c7cfaeff840f360fcbe007c;
mem[136] = 144'h020df2a8f328044ef5ad0069f9fe04f5f3c6;
mem[137] = 144'h019ff99af2d6058efe71f432f27ff89e05d6;
mem[138] = 144'h021c09c706fd023ef01cfa260b55fd8609e4;
mem[139] = 144'h0c91fb2dfc88f6d0f8440c77f380fb74fd1c;
mem[140] = 144'h0ca10ed608a700290ea1033b0fb803dcf489;
mem[141] = 144'hf3e50eadfbaaf490fe3e0384fdd30b7ffaa9;
mem[142] = 144'hfff7061207e9fdd80e0bfaa3f47b0fae02bf;
mem[143] = 144'hf7ab0f8df059f6620a500d98f29ef9b4fc3c;
mem[144] = 144'h00b4fa93f6a801dff09e0623f37a090e071c;
mem[145] = 144'h00660a440849081d0fb9093203f60192080c;
mem[146] = 144'hfd210dda09bd0ac40f85f86506e10ce6fe91;
mem[147] = 144'hf3acf767fd3904def73c0c5d0b4ffa45f11d;
mem[148] = 144'hf9b4fcb9031d0c470f5e0723fc45f17502b6;
mem[149] = 144'h0747ff2e0eb4f1840983f7060b88f88d0dfd;
mem[150] = 144'h0d110b21083704c90536067c07adf6d206f1;
mem[151] = 144'h0e23feb7093df339f213f76c0783f27bf51a;
mem[152] = 144'h081c0888fdc806b1f53a052804850e13fd85;
mem[153] = 144'h01eb0e9a085a000901c90df3049e0f9efd10;
mem[154] = 144'hfec90e57f4280c17f35706860213f991f6bf;
mem[155] = 144'hf9eaff37027dfb49008f0ef50014f324fafb;
mem[156] = 144'hfc48fb240c21fa8f06e5f0680e5e0b86f46e;
mem[157] = 144'h0606fe27f540f598f0ba08b0f6f5f13c0ec2;
mem[158] = 144'hfd2f0bf30662f35d081d0bf4f65a00d2093b;
mem[159] = 144'h09fc09ddfb4bf305fd09f4b601fa0401facc;
mem[160] = 144'hf1b2fc3df1fb0d250d80f94d0b390aa2fdbf;
mem[161] = 144'hfacc07a8f0d002670058f37afa2af58b0b47;
mem[162] = 144'hfe2bf0b9f1abf779f72f0626f658fe2d0510;
mem[163] = 144'h080cf33d0811ff0bf776f99f04200991f0e7;
mem[164] = 144'h08c20378f7e0fdebfecbf32a0ee9ff8d0783;
mem[165] = 144'h0f25fd650a62f25b08c403d700c909900b87;
mem[166] = 144'h0657fc63f99af9bcf5d80287f16d0d570396;
mem[167] = 144'h07f102b602920175088e014ffad2071e04b9;
mem[168] = 144'h02d9f59af162f7d30df8f1640483fd7ff758;
mem[169] = 144'hf2200f030bf0f658096ef597059a0c02fc97;
mem[170] = 144'h03b4005df465efa5fffc0d52fe9ffd5bf88b;
mem[171] = 144'hff2af71ff335f576fee403ad083a054dfa71;
mem[172] = 144'h033ef23ff8d3fb84fc70fb3af2c0fcdf0915;
mem[173] = 144'hf8b7053cf139f26c0da00410fcc4f0fc062c;
mem[174] = 144'hfba40ba1f6a0fcf7f0b60857ef6bfd03f9f4;
mem[175] = 144'h02d3047ef0e8fd1407aaf28c0d2801abf556;
mem[176] = 144'hf9b9fe6af571f4810f4a0626fa55f7bf05f6;
mem[177] = 144'hf27ef5f20b4a0d8cfeb60905027efbce0415;
mem[178] = 144'h06f606fb084b0456ffc8097a0d07f776f612;
mem[179] = 144'h0458fd6bf908005508bff4c0f4d30c87f873;
mem[180] = 144'hf57e0c47eff1f9d6f8290162f1e1095002f1;
mem[181] = 144'h01680878fe6d0afcf4def522f4be03dff6cf;
mem[182] = 144'hf32e07f4f98cf5ddf02a0a300061f5d50654;
mem[183] = 144'h0237f0e802bdf4c7f872054efb3b06cefc06;
mem[184] = 144'h0e34fd22f5f4f7b8fe5c0b73f4d007a8053b;
mem[185] = 144'hf9c0092cfb7bf5af0802f5c6084aff2b08be;
mem[186] = 144'h0d8efd5c0ea7f69ffbac0c3c0e070197f695;
mem[187] = 144'h036df5e1f2a8092def83fc2ffe20f42404b4;
mem[188] = 144'hfa99f9ecf38b0a3a0369fa8afb870661fa01;
mem[189] = 144'h063bf8e7f54df4b9f62d00950c2d02630054;
mem[190] = 144'hf311f27601c903bc0033f4f8fac907b5f1fc;
mem[191] = 144'h02b1025c0a0f0d76fd82fb190521f49bf100;
mem[192] = 144'h086b0403083e0619f57bf05df29bf226f114;
mem[193] = 144'hf4ea0e6f08e4047c06fdffcffe2404f308e5;
mem[194] = 144'h005afa8a0a26f6590ae3fe790e300be0f7fa;
mem[195] = 144'hf7a4f46601bff479fa3b0e7809ff03b8fa19;
mem[196] = 144'hf921fcd70242f90bf35d02d3fde208c8fcc1;
mem[197] = 144'hffe5fc82fbf10774027ef3b40506fb1cfb10;
mem[198] = 144'hf27cf75dfe25f900f14109e80c5b013f0fb5;
mem[199] = 144'hf6f4fc940684f103085100eefa91fe37f4c3;
mem[200] = 144'h036c0ec2066dfa0ffe3df2b9f5a905cefe0c;
mem[201] = 144'hffbbf9cf0ee6f3d4fac90042f9a3f6b6f220;
mem[202] = 144'hf14a0e8108fdf22af055f4e3075ffeedf7fb;
mem[203] = 144'h090c00b0f59e066b09580a82faebf76bfae0;
mem[204] = 144'h0c8bf8a8f93af3a8f2fafe060f520406f4c5;
mem[205] = 144'h053c0692f0a70c7309b9f1c2f96efa23f306;
mem[206] = 144'h09a4f57904a7f06efae60e9af3c3ff7bf43b;
mem[207] = 144'hfa6bf0c20a22ffc1f08d08a0fd5cf740f96b;
mem[208] = 144'h0eb00f9d0565075d0ebc02b5fd6ff8210c3a;
mem[209] = 144'h049ef394042f0876f95bfde6f099f6bcf1e3;
mem[210] = 144'h08daf7aef1e00e77fbda0cc604a0f7e4f307;
mem[211] = 144'hfb69050702d0070c0d8af793fa95f7a7fbf8;
mem[212] = 144'hf1b8f382f118ffae0abf082dfc67068405b4;
mem[213] = 144'h0b0ffc540db705f8fc7b03ee029505cbfbf2;
mem[214] = 144'h0cc107ad07c3f15cf999f0c3f0050656013a;
mem[215] = 144'hf586046af16406aeef83fb8c06d30d1a0531;
mem[216] = 144'hf2c9f7d1fef7f675f9e503d6025607480af6;
mem[217] = 144'h0c40f6daf6d4f2a50680f8adf30f01c1f4f9;
mem[218] = 144'hf45a097df428008409f6f7cf043e082bf5dc;
mem[219] = 144'h0b7bf7ee016f0a57fd1cefcf0aee014feff1;
mem[220] = 144'h0b5df5b0f36dfa08f9aa05bd09d4fafd002c;
mem[221] = 144'h09dbf9c307200820f03efcfdf4dafabdf03b;
mem[222] = 144'hf2e4fd80f1030c490325f10701bc0eea018d;
mem[223] = 144'hf4c6efc2f3b5f86c0142f39d085f0e9dfdd7;
mem[224] = 144'hfd0cf6a3016401f9f79901a8f7b5f72cf067;
mem[225] = 144'h0b77f041ff8bf08b0d430418f0aef136f083;
mem[226] = 144'h06d9ffdbff38013a01bfefb508250649fe53;
mem[227] = 144'hfe91f297f672f7d00067f902fb6af2ccf593;
mem[228] = 144'hf9890acf03a8f294f930f993f50805fff086;
mem[229] = 144'hf941f5cf0c820f5503da00d2f8f1f65206e9;
mem[230] = 144'h0251f1e5fbea047d054f009cf3e2f06af785;
mem[231] = 144'hf6bdf7ef0d02010bf48002cef553f6960b45;
mem[232] = 144'h0052f532f5b3f5b10318eeac0cfdf42cf5f0;
mem[233] = 144'hfffef157faeb07d4f14f06b9fda107d608de;
mem[234] = 144'hf9a0f0ca0940ef26f8c6f6a5f5ae09570e30;
mem[235] = 144'hf1180caef7fdfa35fc6601cafb4efcd5fadd;
mem[236] = 144'hf7f1eed90ecff03b067cef780e8d0da4099e;
mem[237] = 144'hf60af849fd30fb1df66ff2f5f96607050877;
mem[238] = 144'hef28f2ec0e8d0ac10c6407d3ff28fe390ad9;
mem[239] = 144'h0d480782ffe903c7feb9f0840b8d06d70c27;
mem[240] = 144'h042cfed90e570589f3a4047603baf44102cb;
mem[241] = 144'hf25bfc810af9fa8b02a60341f212069b0aae;
mem[242] = 144'hfc8bfd8d04080d44f2a3fc7b030b0eb9f20a;
mem[243] = 144'hf5edf758fdf804480c3bf5160c56f59b01d2;
mem[244] = 144'h0ae70896f4800be1064e0a8af5650de2034f;
mem[245] = 144'hf1a30b00f3d80f6cf709fc790f800525f56f;
mem[246] = 144'hfdfafc8f078cfc9e014bfaddff8c0e0dfe92;
mem[247] = 144'hf4510f35f39104eff4cb037bf3aaf287085f;
mem[248] = 144'hf972fa8cf0130923f06d0ccb0292fe60f831;
mem[249] = 144'hf7bd015b0f90072cf5760c6f0c01f30d01bd;
mem[250] = 144'h09b9fd6a091bfa0ff505ffdd021f01140eb1;
mem[251] = 144'h0bc7027604bff4aa0b31011f0a95fa0c0068;
mem[252] = 144'h002dfe71f14b07600cb905f50bcffd1f0d69;
mem[253] = 144'h080cf37e0ffb0830f7980768f23af3acfe53;
mem[254] = 144'h0243f8c6fa9b009bfc4b041c0e05f3170a99;
mem[255] = 144'hf91dfaa3f29008c3fe57f8e708cd0f160868;
mem[256] = 144'hfa4e0edf04b200d30e14fceb0345f2aa05b9;
mem[257] = 144'hf9f103e4fdf0f8cb0a2ff5c504520ba0ff0f;
mem[258] = 144'hf6010e73f93d0cb80ca907c7fac90bc604fb;
mem[259] = 144'h0dabf2f7fc9209ccfb51044df77902eff4a8;
mem[260] = 144'h04fdf8ac01e50ade033cffb005aaf4090691;
mem[261] = 144'h00430ab4002404abfcaefe06fb8bf0a40ce8;
mem[262] = 144'hf54e05460384062eef25f421f6260a8e07da;
mem[263] = 144'hf9dbf364f76c0f1502bff2bc0dfd0bef0f63;
mem[264] = 144'hfdc1fc480978efdd0c3af765f8eaf329f39c;
mem[265] = 144'hfe060c46f33f090df4fefa54efe70e3bf0f5;
mem[266] = 144'hf08e029b005d030d04fcff390d41020902eb;
mem[267] = 144'h0e2cf6eb0505ff17ff29027dfab3fd4c08c6;
mem[268] = 144'h049df820fd19060c07be0ca2fe62f2310777;
mem[269] = 144'hf58400070dfc05770a68f21bf3130a010dfd;
mem[270] = 144'h0666fe62f4dff1fb0bfd02acefe6ff75f737;
mem[271] = 144'h03e4f6230ad4f53f03fef183fdf3fc5e090b;
mem[272] = 144'h0fbf0d490e170cf0f7c5f73bfdcb0202fe8b;
mem[273] = 144'h0f58fd9ffa5c0848f18df4c1f233f93ff5a9;
mem[274] = 144'h08f60f13fb1bf90e0aa9ee68faa4f645feb9;
mem[275] = 144'hf815f9be0185034ef79b097a09760919f4e8;
mem[276] = 144'h0fd00a3c0d4af567f7910a9a0010071ef993;
mem[277] = 144'h0e630a41fc0efcdb079b0bd6f44ef4120162;
mem[278] = 144'h009cf602f532f8b0f50afa4f0e29f86cf45f;
mem[279] = 144'hfd3d0e62fcdffd820df1f867f19c051ff8f8;
mem[280] = 144'h014af11df2effcf4fd9efb9909aa04def58d;
mem[281] = 144'h089cfc18f2bbfed5f98aefb4f63bf8ecf353;
mem[282] = 144'h0f4d0b71f6da0f34053810710ba90dd4f32f;
mem[283] = 144'hff68efb005cef5ff01aff4acf823ff5304f5;
mem[284] = 144'h08fcf2550de1ffb3046e046f0b9a0ec40130;
mem[285] = 144'hf2f1f903f266fe2b0049f4cb07c4fc93f24f;
mem[286] = 144'hfd04f2c6fa08fcac0462082807b8f8c50f39;
mem[287] = 144'hf0d507e4feadf0ba0d85071b0a5ff602008f;
mem[288] = 144'hfcd700930e4af450052403dfff4ef881fab9;
mem[289] = 144'h0dc804fcf44c07e50a81faf2f715031cf50d;
mem[290] = 144'h00390f34f48bfa62fd7bf60dfda10b190913;
mem[291] = 144'hf580f356fcb70ea1ff0d0aba072ef75303d0;
mem[292] = 144'hfae1f9baf9b80ea7009e0daff35bf706f85c;
mem[293] = 144'hf6f9072e0e100ca60b4803f302d20c1bf958;
mem[294] = 144'hf47af067ff820b560587049c077c064c08b2;
mem[295] = 144'h0a1dfebbff7001df01a6f6e6028309f40999;
mem[296] = 144'h09c3efa5fa52fd4af7b20ddbf98d055ffdd6;
mem[297] = 144'hf26403f4fe1309bff51506430f06095af62a;
mem[298] = 144'h0551f49c0a8cf3ab08290a2d0a65062df9cb;
mem[299] = 144'h01160220011503bcef47018f05e90d02f455;
mem[300] = 144'h07b2fdf20a1305250879f05aff2bf8360e1e;
mem[301] = 144'h09c9031005cf092009c7006c049e0eecf9b1;
mem[302] = 144'h0d8b0182f5c0f449ef62ffb7efbbf57309eb;
mem[303] = 144'hf045f473fbef0861fe39fe0af26306e2f8e9;
mem[304] = 144'hf69002e5f7d70f00ff0403150bd805e7f71f;
mem[305] = 144'hf6da05fa094bffc3040cf09300340739f742;
mem[306] = 144'h0b7208d309e0026e0a6cf60c08e2023d07f0;
mem[307] = 144'hf174037c069df0d7fb90fee70112f5d9fe87;
mem[308] = 144'h0776038ef7b40d990d96f1b4f8eaf29b00d3;
mem[309] = 144'h013400b6fb7bf53301b9f632f32b0892f470;
mem[310] = 144'h05cf060706bbf829f5e005f3ff09035efe71;
mem[311] = 144'h009b0df4f0a7f860ffacfc54f347ff4bfec0;
mem[312] = 144'h05eceff1f67bf369fb7ffa9906c30b5f05f1;
mem[313] = 144'h030a06300b2d04cd062cff880ce601bd0fae;
mem[314] = 144'hff45f102fe6df906fbec0c07042a0bc104fe;
mem[315] = 144'hf44e079ef815f2fa0551f3a2085ef652fdaa;
mem[316] = 144'hfce60f4a04d2f08afa650417fd2a0b0bffbf;
mem[317] = 144'hff430886050dfaf7f50904daf22a07e5f6b9;
mem[318] = 144'hff42f0b6f7a00e9807e3069cfb55f9fe0aa6;
mem[319] = 144'h0c01fcd004170983f5cbfed8040b090ff616;
mem[320] = 144'h029afd2b07ecf441f376f0b30bbcf9e000d6;
mem[321] = 144'hf16effe2fa700f5bf8e8feac0fa2fb1b0e2e;
mem[322] = 144'h0542f922f8380347f9f3f8e7fe53fed4fd6b;
mem[323] = 144'hf18bf035f342003ff8cc0f0108320f80fcec;
mem[324] = 144'h08590b32f93cf70e0a9cf120f6ad0f670b41;
mem[325] = 144'h01060841f68af1dff9a6f2390bfdf613fb9e;
mem[326] = 144'hfa87039c019bf115fe1dfde40efa000c04dc;
mem[327] = 144'h0606fa970fb4efa80b800be0f49700920cf4;
mem[328] = 144'h0d4a0b12f24e090709070388f58afbe3f273;
mem[329] = 144'hf847fa92f1000be205c7fb7900240e83f60c;
mem[330] = 144'hfc2ff2f10756f25c099006a3f2b6099b0d3e;
mem[331] = 144'h0d9aefeffecaf5bbf582045af086f2f90540;
mem[332] = 144'h018cf5c0f5090cdbf10dfe6c0a4df36d078c;
mem[333] = 144'h0572064500b90c91fc7f051a03eb03f60250;
mem[334] = 144'hf34708faf21ffb810e6ef21dfa05f3290f2c;
mem[335] = 144'h0af50bb5fa7df954fc22ffa6f74cf7990b43;
mem[336] = 144'hf734f9b106a20437fcb6fae50a870ea20b6a;
mem[337] = 144'h0c29f846fb5407e4f254fbf2f915fac107bc;
mem[338] = 144'h04a2f32a02cdfd92f727f6700813ff1e0de0;
mem[339] = 144'h0d3afebc0b32077ef857f74af646f4de06ea;
mem[340] = 144'hf46e0de8f45cf8800a06f643072cfb62027e;
mem[341] = 144'h0342feac07be081c0c42f973fd9100fcf812;
mem[342] = 144'h06b70b1c0fd1f5870a9e03bd0abff5750df1;
mem[343] = 144'h023500400d6c07aef12df96d0481fb49f5a8;
mem[344] = 144'h065909c90666fcf4083afd33f758f908f1e7;
mem[345] = 144'h04880428f02affd30bde06370c41092c0828;
mem[346] = 144'h0df10ddbf03af05bf5a0faa6078006effd7e;
mem[347] = 144'hf239f682f704fa5405e2f98806550d31081f;
mem[348] = 144'hfac7f8e7f7b4f5af0a24fef50ed905ac0335;
mem[349] = 144'hfc26f9f40981f303fedf0284fc22036bf851;
mem[350] = 144'hf8510592fb9d095e057b068bf2da0a1ff05a;
mem[351] = 144'h0c3dff13028df631f7650c90f002f542fb3e;
mem[352] = 144'hfeed0bd6f377f394f6eef723043809df0f3f;
mem[353] = 144'hfc0e0ef9fa8405bf0bd9f799fbe1fafdf471;
mem[354] = 144'h0c56068b0859fce20c78f02e0c5efe52007a;
mem[355] = 144'hfa63f4450dbcf5b3f58a070200650c39f995;
mem[356] = 144'hfbb1fd72f9770646f321fde502dff449f826;
mem[357] = 144'h02a80f23022c098c04fd0cb3f866fafc044b;
mem[358] = 144'h0cb803fb0c460f71f8def70601ee0595013e;
mem[359] = 144'hf12fff8f0ae108a2090ff92af06e0f8ff080;
mem[360] = 144'hf9670a49fdbe0770f4af087f01b1f8d20938;
mem[361] = 144'hf726f59708ddfb4d051a0948f6a4fe9f0d15;
mem[362] = 144'h08dff88af868f1a609fffa6cfa5af8f8f9a2;
mem[363] = 144'hf06a0b23fa07f7cd0c6f0259fe3f0cb8eff8;
mem[364] = 144'h0bbaf113f3590439fe42009f0401f5760a79;
mem[365] = 144'h06050c900a62fbfe0361fd310b7f03edf030;
mem[366] = 144'h0446fa780413f346fe2702ca0daefeb90212;
mem[367] = 144'hf9c1fb1a0961f57bf7e3f919ffb700bc0754;
mem[368] = 144'h041bf47cf3db084801d50c32f73df649023b;
mem[369] = 144'hf779f9af03a20e24f8b9fc0af8d0f56b0d0d;
mem[370] = 144'hf404058e006e0d260bbb05da0e59fa3d03e7;
mem[371] = 144'hf7c1f55efafdfa5e02750205f2befcc10b6f;
mem[372] = 144'h07f407b4fad603a2fcf6f1eb0a41fa76f7dc;
mem[373] = 144'hf69707ec08f2fb78f65ffba90462f6c107a4;
mem[374] = 144'h0f8bf03df435f7a7f486fcd5f9fcf80df061;
mem[375] = 144'h09d4096b08f30cf60792029afed1fd1ef864;
mem[376] = 144'h05dc02d80f94060cffc3071d02c1f6ab0654;
mem[377] = 144'hff6cf0a60832f7a2ff62eff305bc0d11f449;
mem[378] = 144'hf396f38a08480e52efffff09feab01f509a1;
mem[379] = 144'hf146f273f934fff10a42098cff45f23af4bc;
mem[380] = 144'h002efe260cbafc2b0f3d097ff5ed0def093a;
mem[381] = 144'hf5280e24091f01c70da80c93f5e2fe02f6e7;
mem[382] = 144'h0857f7fe01080708fbf0fe41040105080f30;
mem[383] = 144'hfba405bffb9df26f052cf3190e98f8b009e9;
mem[384] = 144'h0f0d06b10b27f4f30c5408c702c4034ef9e8;
mem[385] = 144'hf00cf413f826f52706aa08f3f83c0f1ef94e;
mem[386] = 144'hefcc08faf9eb0c2af133f478feb309eb04c3;
mem[387] = 144'hf0f9f39d090ef4720f710408f81bf85af347;
mem[388] = 144'h04b5f288fa26f73cf5f808b5fcc4f6e9060a;
mem[389] = 144'h056dffe30548f15af1c2f9c5f4280944f30f;
mem[390] = 144'h06d40c020071f1f1f1790f2d0dd3f46dfca0;
mem[391] = 144'hf10ef0c5081fffd60a54f5cd061c0b80f0e5;
mem[392] = 144'hff830902ffeaf1ce07fb050dfa7bfe69f073;
mem[393] = 144'h018f06fdfe28fe6206150b2f0bc8f098fb6c;
mem[394] = 144'hf9f10cd50da008150574fa08fd0c0c460e9b;
mem[395] = 144'hfa240bf0fe90fcd2f7c5f8c4071607040e36;
mem[396] = 144'hff6c0d2e0d3b0d52f1ecfded03f300b9f996;
mem[397] = 144'h0314f16d0626fccff00508710f07f38d007f;
mem[398] = 144'hff49fc9efc1d0676f5c6f5dbf3f50ecc0eb9;
mem[399] = 144'h05ab01f0f61409bff2ba0da7faa50a3ff31b;
mem[400] = 144'h0c2bfe8f057c034ff044f26bfffcfd9e0a31;
mem[401] = 144'h024d01bd042900de08880c4ef71106ecfeb2;
mem[402] = 144'hfbe9f8b90644f4df04290f5202e10d9101fa;
mem[403] = 144'h0fcd08920be00dee0a830c1bfd13fbc7f25c;
mem[404] = 144'h0a4c06b909a6f770fc500245f98afe1ff42b;
mem[405] = 144'h0600fd25f2aa06b508d20439fd0903a8ff92;
mem[406] = 144'hf51ff40402bbf43cf451f661fc3f00b2f24e;
mem[407] = 144'h00390194fbd601e80474f4a3f1660cbff647;
mem[408] = 144'hf0430c2df0bfff4e041702d2f902f4710faa;
mem[409] = 144'hf7cc0254f12206560be9f30efdcbfa270950;
mem[410] = 144'hf9f70654f05a0d79fbdcfeb20a660ed0f619;
mem[411] = 144'hf9cff029f23b0db606650f74fc8cf73df323;
mem[412] = 144'hfb22fde9f9550de7006103e6f36df7edf211;
mem[413] = 144'h0761f5470d17f76e0428f185002e0cd1fa89;
mem[414] = 144'h08a10590f771facbf38ef70cfb34f235f324;
mem[415] = 144'h02460dcef92ef1abf60af7c5fa07f34cfe0c;
mem[416] = 144'hf1e90787f86101a8fc9cfd6b0a17fb8ff5a2;
mem[417] = 144'h0ae9f3def9db0bbc08e4f4640937f2eefb3e;
mem[418] = 144'h05c40e30f602f906f3f109e9fe4107950a0b;
mem[419] = 144'h0730f036065f0f94f9230c2b03daf7820c9c;
mem[420] = 144'h0f7f0365fea5f260f8c2f24d0fa80f2404e8;
mem[421] = 144'hf2780cc90927ff90f0eafc330bccfe0ffec8;
mem[422] = 144'hf03d06cbf2e2054c068af507f4b9f5cbf6f5;
mem[423] = 144'hf9180a3ef84ef449fdce06af026b0753f8ef;
mem[424] = 144'h0de80b70f71100b9f1a502da01a6fb4afd23;
mem[425] = 144'h0c65fc5d0828f1a500fafbe5fb26f3e7f716;
mem[426] = 144'hf942fd7ef4dbf0220beef9fdf9abf2d8f780;
mem[427] = 144'hfba6f6b7065e099b0e470376f94306a60c92;
mem[428] = 144'hf7e4f699f1a6f7020bc6064f0d26f9240f3f;
mem[429] = 144'h0edbf318035909f4084b03d40c2dfdbff7e3;
mem[430] = 144'hff4cfe49060300b6fa2fff76ff3af866f626;
mem[431] = 144'h0964fe000724078b08fe01a8fbaff5ef0e8d;
mem[432] = 144'hf99ffc0bf96a0e3aefeff3dbf38afaf901c3;
mem[433] = 144'hf62cf58bf6790e64f3faf492f27803f2f3b7;
mem[434] = 144'hf235f1950d38f3e0fdda0dc7f96af5e50a17;
mem[435] = 144'h0acdfbf5f025083cf73408b4fc06f9390563;
mem[436] = 144'hf732009c06d1f402fff3f00efb0ff52cf168;
mem[437] = 144'hf373086800b10034f870024af3b5fcc50c2a;
mem[438] = 144'hfab8f5f4f2e9f5350b95f872f5d2f3e4f641;
mem[439] = 144'hffc605680410f30f07c2fa760ea109a90307;
mem[440] = 144'hff9af462ff8ef69a06b9f272fe580030033f;
mem[441] = 144'hfa2bfd7ffc2efe24f36bf509f198f05a06bd;
mem[442] = 144'h0e6f0f0d00b9f572f70b02ce095ef2ac010d;
mem[443] = 144'hf4fefa56fff6faf2fd01f856ee9a0380ef3a;
mem[444] = 144'hf44bf17aef6c030ffa52fc42f739f20609f5;
mem[445] = 144'hff33faaef8aa011b071ff9870aa6f313fbfe;
mem[446] = 144'hfacaf485f4e0017aff6d09f9f049f18afdae;
mem[447] = 144'hf947f947fbf8037e0350f60207a702170b91;
mem[448] = 144'hf540fd080f590c7008a205c30b4c041bf6f8;
mem[449] = 144'hfead0481fb78f680f539f86ef381fe4303cf;
mem[450] = 144'hf0c3fbb00c5c02ea0abb0466f32c0885fa2b;
mem[451] = 144'hf211f0360c13f9d2fe9003f1f8faf39ffc98;
mem[452] = 144'hf5adf342fee10f7c065a01700765fba9fe35;
mem[453] = 144'hf743fbf80d670b13fef401010a120bde041a;
mem[454] = 144'h0c790f0806da01030b6f0e4b0795f4dbfaa4;
mem[455] = 144'hf4f3f2ec006ff842038d03fe003105bb0b72;
mem[456] = 144'h0b720592f315f0e7030b0e2a0396f483f77c;
mem[457] = 144'h0b2d0ef508290aa5f3d7f0e80f21f8eff41a;
mem[458] = 144'hfbee0924f36d0a35f992fd77fbb509e20cda;
mem[459] = 144'h0bb4f1500b210f5cfa2009b5fc0c08cafc9a;
mem[460] = 144'h0720f8d60efafbc90600ffba071809dc0cad;
mem[461] = 144'h079d0f0100a5f2da0d0af7fbfedaf1fafde5;
mem[462] = 144'hf6c3f590f1d7f080fc85f2f00f6ef0c802f2;
mem[463] = 144'hfed8054cfbccf9d4067407a6f18bfcb30ae6;
mem[464] = 144'h019f00dff8ec06db05c70f7803e608530545;
mem[465] = 144'h0c23f4440067f41efc47f8ee0db10c88036f;
mem[466] = 144'hff580587fccef470f01efd6b004904f208ba;
mem[467] = 144'h0e63fff90929014a002305b4f4c00704014b;
mem[468] = 144'hf49cf7d308780738fcc00af1f19e0a0d0266;
mem[469] = 144'h069df9fbfd68f517fbd400fe07a40ec009d7;
mem[470] = 144'hf9f7efa6fb02fdb4fdc3065708c5ff450d41;
mem[471] = 144'hf33c0487fc14fa86002bfc05fea600290a06;
mem[472] = 144'h08960bd1f707081df9fbf2820ef8f205f7ad;
mem[473] = 144'h07cef42f07f4071c0306f0d6f784043d01ad;
mem[474] = 144'h0ed105500a540e14fadcf0f2f88602b9fe98;
mem[475] = 144'hf376f305f549f63d014f02f3fabef4a70275;
mem[476] = 144'h097b03ec0cb20a410796f07b0a66ffe5f88f;
mem[477] = 144'h059607a7f5ccf311fa0af89b04c2f37d092a;
mem[478] = 144'hf02bfab5f5a00b0b0caa03d7f9c3f9c4f514;
mem[479] = 144'hfabef6c7fe6afff4fada0d010f740a53f3de;
mem[480] = 144'hf1ba0010f894f8f90fbc0fd0fa3a031ef955;
mem[481] = 144'hf0b60b47f7a20ecbf14d00fc0e6bfcd4f99d;
mem[482] = 144'h08f8fe75089a0796f1acfcca045ff77cff7a;
mem[483] = 144'hff890ba6f3090a59069cf2daf041f845fa99;
mem[484] = 144'hf25507a500e2f71f0def0eb402ed08de0d85;
mem[485] = 144'hfe0d06bffac1f705f98df7240b1406d6f070;
mem[486] = 144'h0c86fb94006901e80f29f05afaf402ff09b4;
mem[487] = 144'h09540527f3ec079df23f007dfd92f2c8f877;
mem[488] = 144'hf941f3a605bbf1e5f1a20fd4f29200e4fa90;
mem[489] = 144'h03b60a39f777fc05f5aa09ab0ad40016f7a5;
mem[490] = 144'h0f38f38805ff0e79fc2ef9c4f27f095103b6;
mem[491] = 144'h014606befe890e71fe50ff8b096b0f00fdea;
mem[492] = 144'h0ef5faf4fd4eff58fb710b4002a0042ff7c3;
mem[493] = 144'h09b0f358f73c05be02fef34903ecf7b6f34e;
mem[494] = 144'h0c9900f4f6b7098f0ca2fb3cf0a20599fe53;
mem[495] = 144'h030b079a06ac0ed10337f3f00309f7660f44;
mem[496] = 144'h0b5af7dcf9c4fa46fe4c029e092df82b0b51;
mem[497] = 144'hff2d086d08fff9b2fdbd0cdffd440c390785;
mem[498] = 144'hf7a1fd0cfe53fb02f596ffd2f52c08e7f032;
mem[499] = 144'h0960f2440a890a02f78bf355f4e40a2a0958;
mem[500] = 144'h0737f3a6032e0c7bff8afdf50872f4effdea;
mem[501] = 144'h009b01bc027cf5cafac2f8f3fd73f918f6aa;
mem[502] = 144'hf41504e0040705d805bcf539021e0b87f6a5;
mem[503] = 144'h0cd50f090838f88bf50ef9b1009bfdb7f4aa;
mem[504] = 144'h0c1201ed0b53fb0d0aa10253075c02f9f0bb;
mem[505] = 144'h049f0957f04fef1ef454fb560a970157eff4;
mem[506] = 144'hf1e707c208b9fa090dfc02a0083c0268f169;
mem[507] = 144'hfc6ef66c0bb8ffa40603f3d700280458fef9;
mem[508] = 144'h087b0761f323f202f0f3faa6f9020cf1fdff;
mem[509] = 144'hf96202d4f7cf0e28fc2103bdff9005370664;
mem[510] = 144'h092eff4204710aecf7f7fe8f08b80c720ce3;
mem[511] = 144'hf9f50ccc0117fbe0f050005e0402014cfb71;
mem[512] = 144'hf140fc27fcbaf1c606690e0b0290ef12fdf0;
mem[513] = 144'hf8caf613066400720886fb46f7dc015408cf;
mem[514] = 144'h0392f703fba2002f0d470b190f1af1b8f8c4;
mem[515] = 144'h05c9f7af098403180c56fafefde203e7f261;
mem[516] = 144'h0d680396f64903d70237f4860ebd01b8fa19;
mem[517] = 144'h0d91f51e07d8f8710cd3fad30f23f60b096a;
mem[518] = 144'hffbbf4e7f11af86bfc02056305df0f5dfb85;
mem[519] = 144'h0ba30b7d0065f6d4f29ef11d07fdfd5ff4f8;
mem[520] = 144'h041c0177fa490994fcf1085a0945079909c0;
mem[521] = 144'hf822f7eff801fa4f0df0021800300f75fedf;
mem[522] = 144'h0416fe9e057af7b0044405c90d3af5d8f55e;
mem[523] = 144'h0ee90b41ef3802050c95fe6d0481f295019b;
mem[524] = 144'hf25efc1507a8f35007c50a61fef9f765fa5c;
mem[525] = 144'h09d3fd66fd32fe8ffd7cf51bfd12fbcafffb;
mem[526] = 144'h0a540d9efa62054607fdf314f14801690fb8;
mem[527] = 144'hf35f03fd0dfbfc36ffbe0cfef10401baefef;
mem[528] = 144'h0c0c0facf7a1054c0530f4520b3c00c0f0b6;
mem[529] = 144'hfddb0374f1e608b30bdaf38cf2cc0afa0d9c;
mem[530] = 144'hf92f08fb0628f5e3feecff1c06f0fdcf08e6;
mem[531] = 144'h0a7cf62df8020e1804330fb10acf00d2f51b;
mem[532] = 144'h037df2d50efefc35feeaf09f054e00bb0f8f;
mem[533] = 144'h08770822fc7209def14405f4f16d08a10aac;
mem[534] = 144'hf97df0fd05900e2300c5007a001cf373f355;
mem[535] = 144'hfb56f5250ee502d70569f82ef7f00e3af2bb;
mem[536] = 144'hf5a6f8400974fbb3f843f343feaaf49df03c;
mem[537] = 144'h0e56f17ff7b5052f00a0f9bbfd02f0a2009f;
mem[538] = 144'hf6f0f4a1f933fb8ef5d4f61500de0411f586;
mem[539] = 144'hfb2207d9ef88efb902dff248f96d0afc01a9;
mem[540] = 144'hfcce02b90bf6f204fbab0d22feb606edf2e1;
mem[541] = 144'hf8eff6a9fcf0077c0abaf05903860f0304fa;
mem[542] = 144'hf5da01040495f63ef02c083c0203f6690f6c;
mem[543] = 144'hf879f4d00a30fef6f0aa02e5045bfc80f963;
mem[544] = 144'hf63e093ff594fedaf1950997efa10d1a0301;
mem[545] = 144'h0b6507b107210117fc3b09310426fa3afdbb;
mem[546] = 144'h073a0e68050ef51201f0f292f93408eff574;
mem[547] = 144'h0cf50ff3f6de0dd1f27af6f8f8130b500e21;
mem[548] = 144'h0d3ffcc10a22f1f7fd03045a092df3e5005a;
mem[549] = 144'h08c5f31af8f6093b0d4df564099a0c1b0ec3;
mem[550] = 144'h05a10063f9fbfdbff44702c7fdc3f3810373;
mem[551] = 144'h0dfcffa1fb11f8c80a9bf5adf9f202cb05ca;
mem[552] = 144'h0168ff050659f9090675fc870d8609cc0350;
mem[553] = 144'hf7b6f8a5f0ad043708a3ff4b0c8405fff5a5;
mem[554] = 144'hfa4d0290f7bc0a5bfba00362fdc102a7fa83;
mem[555] = 144'h0abef3b00d58f95b04f6f554f4c5fc7cf577;
mem[556] = 144'h0a340e330eb0004bf2b705d20b21018008cc;
mem[557] = 144'hfafbfa850f9cf01e0e7bfe81064e04b10336;
mem[558] = 144'h083105cc05d2f3bd066f025e06b3f45601fd;
mem[559] = 144'hf1fe0721087f00c9efb8fcb3043bf8340c3d;
mem[560] = 144'h03550e6c0ea304650bf2fc4d0bce0ea30103;
mem[561] = 144'h0fe407def1cc06e90b0df949fd5af97d0a8c;
mem[562] = 144'h0d95f8e6079b01ff063e0075070404880515;
mem[563] = 144'h0f0f0ebbf8360a9df910faa10746fda50e46;
mem[564] = 144'h0ee60e140d6209b20c680d45f57303fdf0c1;
mem[565] = 144'hfb92f42605c1062dfa55fd640d59ffcc0a82;
mem[566] = 144'hfef906e0f941fdcf0a410e3af99504ccf874;
mem[567] = 144'h040d09240b4d04bf09fd011809e5060f0fb3;
mem[568] = 144'hf093f73bfb4cfaa4044bfd9b02810ce0f62f;
mem[569] = 144'h019b0ea5070b08a9f6d9f28af72304b7f218;
mem[570] = 144'h09d806e7003d0613036a03cf080c0cae0267;
mem[571] = 144'h0cd0efe808c0f233fb6a0876fc07f136f41a;
mem[572] = 144'h0c17fcd2fdb3f0270537f4f90c1c0b0a0937;
mem[573] = 144'h0a3601a0fc46f7b20681fa89f89b0d75fa19;
mem[574] = 144'h083a0323f1a3fa850d160e07027efac100f6;
mem[575] = 144'hfb6107d5f2c50fcbf787033ffea7f59d03c8;
mem[576] = 144'hfd8dfa790305fcc6f6a3005807270faefa6f;
mem[577] = 144'h0c430436f3740b9ef56e07e9f221086f01be;
mem[578] = 144'hef5c0cf6fe0f02b50d9bf3a108b703edfcf3;
mem[579] = 144'h08420f5bff820b1e0122074d027bf7a40cb4;
mem[580] = 144'h07650deef18b00ccfb520e4ff555fdb10098;
mem[581] = 144'hfd41fc6004deffeb0b09f3ca064cf02b04ff;
mem[582] = 144'h0e81fede06440b400bb1fe5aefbd027d0731;
mem[583] = 144'hfbacf869f3c30434f235f33afc49f52803a9;
mem[584] = 144'hf4f2073a0017f2a201e7f09308d30fb40aa1;
mem[585] = 144'hf41af3baf32e0a59fb430c3c066ff9f5048f;
mem[586] = 144'hf419f685f17bfc78efe7fe3908960cb503b8;
mem[587] = 144'h0762f837f2f4fe99014f064603a40a2d0941;
mem[588] = 144'h048cf4da07b302c80cfb0872007004fc055f;
mem[589] = 144'hf8c9f59502b80a880d09fe2e0ce103e3004d;
mem[590] = 144'hfb32f94df872f96a0d650d3f069206660f59;
mem[591] = 144'hef59f98df0dafada00f505c1fdf4fdc1fb12;
mem[592] = 144'hf75403d5fb9f0070fd63f2220239ff1a0dba;
mem[593] = 144'h09ab07670388f61f0a54fa3df57ff115f2ca;
mem[594] = 144'h0e840cb30ae7ffd0eff1076bfb3b02c7060e;
mem[595] = 144'h09e7fc8a07680beffdd004a2f8860f670f32;
mem[596] = 144'h025e0b1ffb4305fdfe36f14208090422fa88;
mem[597] = 144'h0278f954fb7fffe700a3f77e084f0a36f72b;
mem[598] = 144'heffe02ddfed0062cf562059cff72f3e5fb1e;
mem[599] = 144'h0f4cfa350ce7029b0a39f95407c300f2f189;
mem[600] = 144'h06c0016905dbf5ad096dfde6f1d8fb3bfa15;
mem[601] = 144'h02baf56303a10819087ef4b40a97eff2f823;
mem[602] = 144'h0eec0318006ef692efb0f483eee307d1f25f;
mem[603] = 144'hfb43095708200389f714fbc00dde0b93090f;
mem[604] = 144'hfd2bfe8ef681f562fd30fa460a93fdb10b20;
mem[605] = 144'hf5520518f07c05050494eff4015e09c9fd85;
mem[606] = 144'h07effee4089b0334f97206de05be0ab6004b;
mem[607] = 144'hf27b0273f1f7047e0ceafe620969fdd4f272;
mem[608] = 144'h0c9000760c30f652065affb6f31a04360a66;
mem[609] = 144'h0d480f8e0b510e060215feb80dea0ef0f036;
mem[610] = 144'h0cfd017ff643f16a0e35fb61fea806e4f3c7;
mem[611] = 144'hf680f7d8f6c2f3f8f5ecf27c076b0b6304db;
mem[612] = 144'h062700e8f854f706f7800a3200d2fb2a042a;
mem[613] = 144'hf9ccfc9df0cd088b02cd03fffc00ffe8fdc0;
mem[614] = 144'h01030753fd920798fc2205da044102da07ea;
mem[615] = 144'hfb4bfc3c0d4502d104a7f86308a7064d084f;
mem[616] = 144'h0908f3e1fbc6f7eff2f802baf51efdd80674;
mem[617] = 144'hf778f332fd0ffe30f15df311024e09610950;
mem[618] = 144'hf1b7f2970c6307deff7e0531f016f77a092d;
mem[619] = 144'h0df4fa6d098604d90f90faeef29b02e8003c;
mem[620] = 144'hfd73f6d7f9310d7bf0860d940a5a024ef695;
mem[621] = 144'hff52f1abf2830ea80da7086e0c9ffdeaffed;
mem[622] = 144'h014ff04ef6d50237f2d0f9170ba605e7071a;
mem[623] = 144'hfb96029c095e006bf1da0e51043ffc63f590;
mem[624] = 144'h089cfc41fd880ed20886fd64ff5b097703e7;
mem[625] = 144'h067d094d03c5f921f72a085eff91f778f7c0;
mem[626] = 144'hfcb8fa80050901f8f17106340a5ff497fbf0;
mem[627] = 144'hf0910a41f3b2095e010f0cc70ab6f9f90a78;
mem[628] = 144'hfab2ff0c0567f803ffa3fb50fc9ffa2c00e7;
mem[629] = 144'hfca501a600870323f0f2fd2af29ff569fbc6;
mem[630] = 144'h033d02b1ff100457fb17f001f4f2091d0d62;
mem[631] = 144'hf8cb0575f8e1fe1ff7fffceff4aef979083c;
mem[632] = 144'hf032f462fccf0a50f7c5097c03bff85006ef;
mem[633] = 144'h053c03140f0dfdf800d3f93f0787ff24fcf8;
mem[634] = 144'h0e4a0a490d9907c2f3fd007ef7faf6ff0359;
mem[635] = 144'hfc10f91efc1cf4d1051e07640734f59df344;
mem[636] = 144'hf554f4e6038108bff817f82ff348fbb104b0;
mem[637] = 144'h0d5fef9b08f9077b0c9b086cf2fe07d80c58;
mem[638] = 144'h083c0152f91cf798f7f5f85df3b6f2990b13;
mem[639] = 144'hfd3e0ee607c9082ff59df435f5f105ac0ab6;
mem[640] = 144'hfa29012001820db4f946f6bd05e3fe870f8f;
mem[641] = 144'h0b4dfdb9f4c00ac4062ff88bfe7efdcbfd52;
mem[642] = 144'hf037f4a101b00d5bf1b808fd0c130270f00e;
mem[643] = 144'h083d0c380150fc7cf942fae10a8609f7f967;
mem[644] = 144'hf86cf826feac0b20fa690da3fcc20ce20783;
mem[645] = 144'h0c14fc0106f10261f30efb360386f6bc0fb0;
mem[646] = 144'hfcb2f684f530f448f5a4f3c1043f0ab5f162;
mem[647] = 144'hf417f81800870afaf029022eff8dfc4e0e7d;
mem[648] = 144'hf67c073cf2b904560429f411f45ff95bf6ac;
mem[649] = 144'hfa2bf831fcfe0f500a11f92dfb84f20c081a;
mem[650] = 144'hf531fc5cf4780b60efcc0b9ff788083af4df;
mem[651] = 144'hf069f63ef899fd5a05e8ffd2f74d096e08a7;
mem[652] = 144'hf69707fc0bb3fa3df375fa98f7e6f7f70486;
mem[653] = 144'h02fd029c01da0ce201d50596f2470d5bf818;
mem[654] = 144'h0f41073b0d6d0bd9f5f60707f5cc0b8bf703;
mem[655] = 144'hf7960d63faa70350f4b0ff990ee704e2f26a;
mem[656] = 144'h0e890247fb6cf7010f3af6580dbff4eff8ea;
mem[657] = 144'hffa6fa85f361f94cfb0c07f00509fce70856;
mem[658] = 144'hf13b0c94f936ffd90cb10c4204080849fb73;
mem[659] = 144'hfc57060c0516007a063c00a7fe58f34bfcfc;
mem[660] = 144'h0c5a004e0c07fa1c01360801f12106e7f4e9;
mem[661] = 144'hf16afff1fa9efd5e009c0968f5f60e2d0585;
mem[662] = 144'h028eefaf018b0a34f9a9fe13f1a4f162ee07;
mem[663] = 144'hf2b0fd3c0e7cfbcb04a50fb0f17ff7e6fd7c;
mem[664] = 144'h03dd01f708810da3079eff6d01c003b30692;
mem[665] = 144'h0b3603670b0808cafdb20dad02def715f86f;
mem[666] = 144'h051b037ef76d0c09f733072a00faf8770d01;
mem[667] = 144'hfbe6fafe04f5045ef97ef7b20949090a0d7f;
mem[668] = 144'h0b2bfb2eff55f9430d2cfcb20ba0f576f30f;
mem[669] = 144'hfb25fa27076f05f507c50150f72802c9fe16;
mem[670] = 144'h059d07e90951056b063c04e105aa0d6df9ba;
mem[671] = 144'hfe6af86e009ef57d0ea2f10f00baf7f00ce1;
mem[672] = 144'hfeb4f03205f70a20ff1108d1f06bfa5e0afc;
mem[673] = 144'hf9b7f11401f6ff30f15c051cf62c0afcf076;
mem[674] = 144'h0891ff0b085003e0f757fab2f3d4081e00e3;
mem[675] = 144'hf7120b65f51df659f05c030ef696f13001ca;
mem[676] = 144'hf8caf5a10781f5b7046800a80511fece07f2;
mem[677] = 144'hfb3ef7e2065af0430e2ffab603b0f2630727;
mem[678] = 144'hf5f0f9890e6cf33a0af20a45f454f2e2ffcd;
mem[679] = 144'hf030f515f72f098ceffdf1e3fde800f4fd70;
mem[680] = 144'h00ad03520799f71201c8f2ef0732f6b207b9;
mem[681] = 144'hf067ff89f25b03eff2a20a99f46dfee609fe;
mem[682] = 144'hf186fff9f95408e406ff0cb0f2a8f4eef124;
mem[683] = 144'hf1e400410983f56a0603efa7efbd0ae7f09f;
mem[684] = 144'hf9ec061afaec0669ff7c02f703c8f25f04b5;
mem[685] = 144'hf4cdfc1cf3aaf09ef834ff65fd62f2f209bb;
mem[686] = 144'hff030844fb5307d0fc6aef8bfa45fdae004e;
mem[687] = 144'hfe41fa10f85505b30b70f4a2f8affab5f1b7;
mem[688] = 144'h08bb02f00c10ff8ffecbf608020ffcc60a9e;
mem[689] = 144'hfc69f0e408fb0d9400a900b6f889f2c00b96;
mem[690] = 144'hf98cf2c0fdebff49fd75f28b0191071cf7c8;
mem[691] = 144'h0ccdf21ffe53f08ffd370a61045703a00e2c;
mem[692] = 144'hfca4f24ff3b100be02d60dd6f532ff3404bd;
mem[693] = 144'hf5c1f6240231f107fa5404620a23034d0a99;
mem[694] = 144'hfa9a09d6f1beff390bcdf2fff80a0ae704b1;
mem[695] = 144'hfe51fcc8064ff47302fbf33f08ab0e1dffc1;
mem[696] = 144'h038af3f7f88e037efeb2f0eafa8f0c20fdee;
mem[697] = 144'hf86c0d66019d0c45fdb8f8df03b2f56ef8a0;
mem[698] = 144'h0f360f09ff85fa9ffb7ef1f9f8ff02d4026c;
mem[699] = 144'h0d41048e0d5c0f85fa29feb500b30997f72e;
mem[700] = 144'h072203e4f7dbf85bf28cfd38f1f1f468f3dc;
mem[701] = 144'h075e03ef0188f2fa0b4af363f4cb00d5feed;
mem[702] = 144'hfb240e6c0b6d02650a7af598076a0bcb0d51;
mem[703] = 144'hfca9f88203b40ae3f1d70183f4590adb09c6;
mem[704] = 144'hf1b5f6e40251f41a0597f835fe360a860341;
mem[705] = 144'hf0d6fb07fa85f1cc048afa20f29f07bcf40b;
mem[706] = 144'h038c01e401a901c5fb8bf0000651f64a04bf;
mem[707] = 144'hf413f84d0515008f09a9040e0538f2e4f771;
mem[708] = 144'hff55f3c8f4daf87cf4d1ffcafa72fd8bf28d;
mem[709] = 144'h05fa054ef7e001ecf639f9000e4e00c4fc1d;
mem[710] = 144'h0699f3d6f940051d05b0f2ef021df554f993;
mem[711] = 144'h0586f9c7f6fef7dd0d5c03b20313fd4bf76f;
mem[712] = 144'hfb2aefe8fd62f73c0589008ef476f4e30920;
mem[713] = 144'hf2d90d310eb8ff690a2d0f0cf6420bc00a82;
mem[714] = 144'hfec60265f64cff6cf3b609a70eeeffcaf7e4;
mem[715] = 144'h0e14048af17df165fc15f2a809ddff3dfc72;
mem[716] = 144'h09a6f723fd600ec4024502c10abf0ad3022d;
mem[717] = 144'h04150366feaefbbc086c0e2cf4c0f96b0ad3;
mem[718] = 144'h0c980f2ff2dafa7d0a6af30bf7e3ff49f0b7;
mem[719] = 144'hfb640804fe55f3440a7b05a507dc0718f654;
mem[720] = 144'h0fadf6b10a50ffe0f202feec0fad05260365;
mem[721] = 144'hf615feedf7040ad0fbf60b98fc42f2e30609;
mem[722] = 144'hf365fde10d070684f5d6fefb05bdf56b08a3;
mem[723] = 144'hf9d80f5a0d1e0707056b01fff515f80df351;
mem[724] = 144'h0f09f796088606fcf3d30cfe03ec071cf72a;
mem[725] = 144'hf9b5f6a2fd4ef63efb99077f0c880dddf4ea;
mem[726] = 144'h058df6ba0696f29c0a63f8ceff77f0cf00af;
mem[727] = 144'hf819fe63fbc6ff16fa6ef342fc6e018dfee3;
mem[728] = 144'h09120ea0f2410ceafa520bc7f00001d2f703;
mem[729] = 144'hfb51f74e04d9f302f66a03a0febff1ae01c6;
mem[730] = 144'h0156f1acf1c5f809030a062a030b094f0d7e;
mem[731] = 144'hf602016802ff0542f0b50333f20b0da0f0da;
mem[732] = 144'hf9e6fbcd00dd0c800172057f00be0a88f112;
mem[733] = 144'h05880f36f664f1fcfffef88e06c4fd21004f;
mem[734] = 144'hf801013efc4900890f2af208f96b0f44f7ea;
mem[735] = 144'hf8e00023fe57f3710bb50df2f559f169f729;
mem[736] = 144'h03d907caf32707e40fb0fadaf532f5c50bdd;
mem[737] = 144'h05d6f90ff960f1690af50262f528019c066e;
mem[738] = 144'hfa090acb08d5fbbdf36409f70490f46af9c7;
mem[739] = 144'h088cf31cf57900b4f170f4cef0360c5effa4;
mem[740] = 144'h00cd0358fc0b009001b8075cfcc80f06f58d;
mem[741] = 144'h0aa5f807fe240089ff9f02c707a106c009f9;
mem[742] = 144'hfd70f95206b8f74cf553f64101fdf662f7ec;
mem[743] = 144'h0b55f90a0cfbf85cf2fcfc19018cf9adf298;
mem[744] = 144'hffe5fdc0f20cf3c1faeaf0b60dcef7c8f3e4;
mem[745] = 144'h062afafe0cbe05ccf14af38b02a90dcbfcb5;
mem[746] = 144'h05d8f008fa6001f8fca2064bf6f90d410965;
mem[747] = 144'h0b8c090c09e5f52707f601810d93f4920b0f;
mem[748] = 144'h06510aa7065b0e62fb080210f92b075dfbdc;
mem[749] = 144'hf4260329f7e4f6c003c4fa2ff4ac05500229;
mem[750] = 144'hf003fedff4c3fcc5f24309d20cc80712fe04;
mem[751] = 144'hfeb10a87fd27f12e05c2f9470a230ea80bc1;
mem[752] = 144'h0e430c970d29020a0ee2f84d08e30910f12f;
mem[753] = 144'hf7f8f4c1031704400f9f03530047045a0979;
mem[754] = 144'h03edf0fdf76b040601a30311f8c305f0f419;
mem[755] = 144'hf36603ff0a0c0b08024300640cca0f13ffee;
mem[756] = 144'hf873fac403780144fc1afbeff0a20f8f0afc;
mem[757] = 144'h0115f62006ba0a26f2a001fdf1b2f642fbf5;
mem[758] = 144'h0575f314eff70dcff3f0f66ff42c0af3f755;
mem[759] = 144'h03150879f23f01ec0b1a0c8dfb9002acf7ad;
mem[760] = 144'hf8240f4f0e0b03cb0202050ff60f04c40adf;
mem[761] = 144'h07b3f87208540c510870f1c203d7feab04f2;
mem[762] = 144'h0f9600b2f1befacef2a5f8b2036601710a97;
mem[763] = 144'h0d02f72f03a0f5630cd2faa403a008abf8b8;
mem[764] = 144'hfab5ff0703660b31fdd6042207da0079fbe5;
mem[765] = 144'h0459f51505d3f88803e902b105e2f834f264;
mem[766] = 144'h012ff80206d8051d0cc4f9f20516f607f647;
mem[767] = 144'h074504de0ed3028bf132fa7dfe230d6c089c;
mem[768] = 144'h0b59f183fd39f47f06970998fb6bfe5a062e;
mem[769] = 144'hf72c0dc3005908e30d8dfcaaf6a009390d18;
mem[770] = 144'h02bef7cd02d0fe41f51402940a73f0a00019;
mem[771] = 144'h01d5fc42fa930d380ec6f02aff8af517f1c1;
mem[772] = 144'h0b1dfbb00c3df04af7fefe37f96d0933f1b7;
mem[773] = 144'hf56604a1fc44ff800794f5c803140f91f334;
mem[774] = 144'h00400115f8d3f9cdf9a4089a02adf2ef01bd;
mem[775] = 144'h0df2fcf10427efec0d000f8f0ae3f18df0bc;
mem[776] = 144'hf859f6f6053efc240a360e7e097508fc02da;
mem[777] = 144'h034304a002cf0097f0220bd7f4620384f724;
mem[778] = 144'h00a3fb4aefd60b4a0034f99a0721f95b069d;
mem[779] = 144'hff550b55032e0b3dffc8f62efafdf5bf094b;
mem[780] = 144'hffd108b8f16af687fca9fe33f0fffd6af705;
mem[781] = 144'hf19509e0f48bf410ef6af8f8f7d7f9db0875;
mem[782] = 144'h04bafbd6fba3f7c5f2f00e68016dfc61fa50;
mem[783] = 144'hfa64f455085800c5f8640300f2cbf4b80e51;
mem[784] = 144'hfff8f247f1670fa9fc6ff864fe730ef6fd23;
mem[785] = 144'hf691fa59f620fdf2f21604c90dc800830d64;
mem[786] = 144'hf4ecff3e03e8f3f30a5602ac0adcfadc015b;
mem[787] = 144'h0209f3cdf097fb6808a4028ff580f500f2fa;
mem[788] = 144'h0314f38c0ef10a9304920e9ef353f139f920;
mem[789] = 144'h0cfcfd92f95e0af7f6e7014bf92bf38df4eb;
mem[790] = 144'h0939f8fafb7a0338f3c5f2b1040afd66fe22;
mem[791] = 144'hfaecff44f56604150d71055e06e90adc0bcb;
mem[792] = 144'hf070f306f332065b0282f22cf375f28ef21c;
mem[793] = 144'hf6150818026fff5a0cfe0ec70569f00ef0d8;
mem[794] = 144'hf6f80e2d0a0ef5ef00f0ff32f4e50725fdeb;
mem[795] = 144'hfe98f461fa01fa69feaefbe80b0df54cf7f8;
mem[796] = 144'h0afb0cf20cad07eeeff5fe89f2f0f20bfb5e;
mem[797] = 144'hf0e6f213f89ffb37ff4d04d4f4aff87afbfa;
mem[798] = 144'hf037fafa093c0cde0de709c0f562f3030440;
mem[799] = 144'h0391004df6f60b46027a0cc3fb81f567fd5d;
mem[800] = 144'hf0bf0c7a0f610900fd0df9020ed6f26dfc23;
mem[801] = 144'h0ad60f310056f9e80d5bf082fd630300f26c;
mem[802] = 144'h03590ce1f96af00905560e960750fff20baf;
mem[803] = 144'h0c2e02580bb7f909fd2b0f9b0e3cfd19f373;
mem[804] = 144'h0a1cfbf108ebf9c909c2f9d50506f7c3f595;
mem[805] = 144'h0be3041bfeabf855f401fe79ff8cf8950209;
mem[806] = 144'h0856f119021dfd99feaaf91d0c42f5dcf54b;
mem[807] = 144'h00c4001304ecfd8cf0abfa5afd200c9b0e52;
mem[808] = 144'hf552fdc70f11f6880090f93f05540b5d067d;
mem[809] = 144'h0a920d5df0a3fd09ff5bfa59f1dbffe10b62;
mem[810] = 144'hfc26f606f7f70028f07802c20891f438f9c6;
mem[811] = 144'hf3f4fbb8f729f0b2ffd7f4adf242fcbc0d77;
mem[812] = 144'hff73fa4e046df16107f7ff050363fb8afd8f;
mem[813] = 144'h0c0ff158fcd5f3a5f91ef3f2f91dfb240409;
mem[814] = 144'hf00a0f3df9780a150ac903d40c38046f0ddc;
mem[815] = 144'h0103fb71f98af7c504e4f81109620d66f997;
mem[816] = 144'heffff93ef0b0fcf4fca4f2c0f602ff9cfc24;
mem[817] = 144'h091f09a20d4ef4bb07fc0b75fbd1f54ffd40;
mem[818] = 144'hf651fb6a04f6f01f004d0d7d05a10b6f01d7;
mem[819] = 144'hf23cfdc80ceefec20f2df79bfd77f4560357;
mem[820] = 144'hf48406f701bcf34cf183f442011bf4c407b7;
mem[821] = 144'hf07f02e1013ef0f7042cf578f82afe57f5bc;
mem[822] = 144'hf9bff58bf482fc0d0325f21f033205040acc;
mem[823] = 144'hf8b4f676051f0ab706e103bcfeb80d48f0e6;
mem[824] = 144'h07660e49f96402acf3a50db5fe3409cb0e03;
mem[825] = 144'hf51801d1027009c808b1ef340d00f3040ad7;
mem[826] = 144'hf27f0a2403980d00002d0ccafff8fc26053a;
mem[827] = 144'hf87002d8fd670e81f3180ab1f899f1e20d08;
mem[828] = 144'hef3e01ba0b6ffe4c0d7b01230c130e170642;
mem[829] = 144'hf4a209a3082fff2f0f0c02e0ffcc0615fcf9;
mem[830] = 144'hf236ff9bf34af48af35301ca0a2ff0940e99;
mem[831] = 144'hf2cbf705fd5cfd560705f13e042df6560a04;
mem[832] = 144'h0da7f7a404e7ffd5fa70f0d2fd18f39bf5b3;
mem[833] = 144'hfc8ef2e4fc1d0755fe290be60098077e0136;
mem[834] = 144'h04fcf04dfdb601d6f8ac0a4b08eb0a900467;
mem[835] = 144'h077704fd04580bc1fdf6001d0a4c0662f9e7;
mem[836] = 144'h0a45f6f5fb3ef76dfe5b01f301baffe203f7;
mem[837] = 144'hfb950998056a0fdff2c3fcc400160097f23a;
mem[838] = 144'h0eb5f0ee0823f6dc07ce0847f2a2fde5fbc6;
mem[839] = 144'hf17d0d2f03c10b110d8bf7b5f248099bf5b3;
mem[840] = 144'hf5fcf76ff1d0fd69f40d0a3bfb12f8e7f731;
mem[841] = 144'hf305f9710adcf04cff2e0c45fd7e0d43ff4c;
mem[842] = 144'hff93f5caf2b9f1cef7f8060d0c1b0458f86d;
mem[843] = 144'hfe79f179fcff08f507d303080c67f4530b2d;
mem[844] = 144'h0b41f45af0e60d5ff9670096067af91df206;
mem[845] = 144'h0bcf0820fbabfb76f6e1f4ac09c1faccf0dc;
mem[846] = 144'hf5a4fbcbfcf3f798fe360adbf412fdc4079d;
mem[847] = 144'hefdbf44af394fe4b02ff07d8faddff35f9f0;
mem[848] = 144'hfeb2f05afb290225fafc0e05f37cf8cb0af1;
mem[849] = 144'h06b20c74f39a0c90fb26f8940eb3097102f9;
mem[850] = 144'h0394f2350aa2f780fc80ef4903da0ac5fc4e;
mem[851] = 144'hf474096b0479031d023ff58efd8bf2250385;
mem[852] = 144'hfdb6fe10f8a50a5407cef533fc4b0279f702;
mem[853] = 144'h0a5bfeda087803fef76c006a0ce8ff0bfdfd;
mem[854] = 144'h01be0cc2f05af4b6fb520d6df5da06a9f538;
mem[855] = 144'h04bd0898070c0178faf80b14f3160dce04cd;
mem[856] = 144'hfe07ff6a092cf342018bf1db0f5bf7790552;
mem[857] = 144'h096cfcddff8b0290ff760a6e01aa00230779;
mem[858] = 144'hf2790104094808990c4ceeee033bf027f3d0;
mem[859] = 144'hfe380c780a9e0d0802d1fe7bf960fd56fb8f;
mem[860] = 144'h02daf429094ff865fb1ffbb0015c0e760ac4;
mem[861] = 144'hfef4ffc601adf3af010cfef1f6610a580be6;
mem[862] = 144'h092b062d0e41f1730a170b6b032bfc9b0190;
mem[863] = 144'h082a007c0643f852f964f8e60ce5029df11b;
mem[864] = 144'hfe590b9bfc2e0333f1f2fd0707f70acc07b4;
mem[865] = 144'hf71705d1f90b0bdbf7330d9dfe6bf192074c;
mem[866] = 144'h08e8fd08f04e05d9f63af172fdecfd11f2fa;
mem[867] = 144'hf562f606036dfa58f0ba06b8fc2a07720c64;
mem[868] = 144'h0914fe5b0d7ffff80862f8aefb610df0027f;
mem[869] = 144'h0e560f0efa8b0eb90f9101350ccc00880c1d;
mem[870] = 144'h019c0115efb6004f0349efbef459056af229;
mem[871] = 144'h0422fcd8f5fd0792f773f8c40e9b04c6f471;
mem[872] = 144'h0940f53bf3fe0539016f052af6ec0b3e0116;
mem[873] = 144'hf5c2fc2c0b09083006c9fc23fd44fe40f984;
mem[874] = 144'hf2410a52fa020729fc53ff720da5087efecf;
mem[875] = 144'h0c1ff0acf4ae000bf0fe0a96054bf72ef8d4;
mem[876] = 144'hfc8bf999f409f39ff7fb0debf424052301ac;
mem[877] = 144'h0363fe58030a0380f630ffa70be00cbe0149;
mem[878] = 144'hfb7cf9630bccef98fd2ffecffdbcf239f60a;
mem[879] = 144'h054206ccf3f9f4f7f13803a9ffa102c1fb88;
mem[880] = 144'h02d606ce0a59f0e904ec0c8b082ffeb400ef;
mem[881] = 144'hfb5202b80da1fa5bfeee048ef093f5adf7f4;
mem[882] = 144'h015000e503bafff1f4d2f87ef6c507610804;
mem[883] = 144'h0a4bf8aaff02f796f6a001f3fd6a0278f0ce;
mem[884] = 144'h09c70427feb4fdc20712fc8c078cff40ff08;
mem[885] = 144'h0f470f2efede0b9bf6eafbc8fc0f0a16f32a;
mem[886] = 144'hf1dc03dff4780e140c54f2c0f83d03b80384;
mem[887] = 144'hfe0505f60d22f33004cfff7501d80c8d02c9;
mem[888] = 144'h040b05dc0fddf158fe75f5340efb0901ff6e;
mem[889] = 144'h0d2cfe4b06900958f750f0500c040ec1fa73;
mem[890] = 144'hfbda059909140559069ef7e809c50715ff53;
mem[891] = 144'hf33008110620ff7ef8adfa820a5c053ff942;
mem[892] = 144'hf2d9efee0eed07090b330a33096f0f2bfcca;
mem[893] = 144'h01c4fc340800f5d4019a0d9bf8af0e0df6bc;
mem[894] = 144'h05a1ff16f26af91df6ae09cafe86058f04a6;
mem[895] = 144'h0b8efddbf31ef0aef568fce9fe98f9c507c7;
mem[896] = 144'hfa72033500aefde004c00e820bb106b501d9;
mem[897] = 144'h0793fcb9f7a107d0f7d80c08f505fd410e7c;
mem[898] = 144'hfcc90a7b070a07bc06e50ae20c96f6acf028;
mem[899] = 144'hf4400219f0ac0cd4069a06980bc1f4d705ba;
mem[900] = 144'h049906300858f800f49f0bd2fe6afbc80083;
mem[901] = 144'h044cfcc70e44fb94ff96f6720d3a0fe3fa22;
mem[902] = 144'hfa9b0d780f1afb8d0dd2038afca706aa0f22;
mem[903] = 144'hfecb0baff4ec03b6fec1ff29f6e1084b0a33;
mem[904] = 144'h0f81017104b4f276f4cafbe8eff7f53b0808;
mem[905] = 144'h06cd0892fb820ca707e3f63bf81ef3b90f42;
mem[906] = 144'h03fb01b302d3044405ad085304850d5909e0;
mem[907] = 144'h0fa7f539fd130a4cf66af29cff170e140c28;
mem[908] = 144'hfd08fe2efbaa09d10245f5f9fbc0f6fb02c9;
mem[909] = 144'hfa27f826fec1f362f5700df2f3d1f0be0abf;
mem[910] = 144'h071ef1140bb8f91df3f303cdff61fa39f3a0;
mem[911] = 144'h0f43f62c0e6908650d51fa7af9fafcadfbde;
mem[912] = 144'h0032f37bf5a00a42fbbb0640f6220614ffb5;
mem[913] = 144'hfb4a089e02e2f102040902f400eaf0fc0203;
mem[914] = 144'hf4dc0833f77a007ff132fd5ef951fb5bffbd;
mem[915] = 144'hfb5c0704f4e5015001e80a67049c0e240e64;
mem[916] = 144'h0555019a0af9fd6b02b00bf5fa7d0c3ff03a;
mem[917] = 144'hfd8a0bd9092cf5a7f3770d84f537f8c60cac;
mem[918] = 144'hffdbf217f09ff7b4074ef45d056609a5f5d3;
mem[919] = 144'hfd96f0d3f211fb79fb2f069d0f4ff56a03eb;
mem[920] = 144'hf940f297f825f784081900f8f56505b3f0d6;
mem[921] = 144'h07c2f519fcf6046a0c14f80a029ff60703f5;
mem[922] = 144'h043ef18cfd53093509daf596f90f0b10018f;
mem[923] = 144'hf40a0aa40176fc00f01809aefa18f92005ba;
mem[924] = 144'h0851016aff4c0baaf0c5f622ff29f5befe5b;
mem[925] = 144'h00edf82f0dd40070034df25bef67efd30cd5;
mem[926] = 144'hfb770af609420b56f44affaaf0800c0bf616;
mem[927] = 144'hefcd06e2f46fff0106c3f2c8f88c0ee6f742;
mem[928] = 144'hf3f50876f496f75a0a34fe1200730434f083;
mem[929] = 144'hf60bf426f219fe720d7a000ef4010b2d098e;
mem[930] = 144'h0c05fc82fadcfd230697080d07bbfff9f506;
mem[931] = 144'h0a800db3f3e1f81707fcf8a8f0810b71f121;
mem[932] = 144'hf7a9fcc80289017ff9a1077c017a07980461;
mem[933] = 144'hf733f63c012906c401a8fddf0171f135fb7b;
mem[934] = 144'hfbc4ffefff320d0f0de2018308610eddfbe4;
mem[935] = 144'hfc82f76a06a0f16cf4e1fde2089fffb80d74;
mem[936] = 144'h0bc9fec3f5b4f8c5fc0d09c8f221f7140425;
mem[937] = 144'hfec0fac100f8f139f2abf82af202060907fb;
mem[938] = 144'hef41f5d704e9fa190ea1efca083cf256fa9a;
mem[939] = 144'h0b310ab5f8cc095e039df9240899f9030339;
mem[940] = 144'hfc690f51ef3af7d1ff79fbe5f937fad003d9;
mem[941] = 144'hf089f3ca0c06f79300160e650c0ffbaa01c3;
mem[942] = 144'heff0fe2508650905f12e044cfb86f53c0964;
mem[943] = 144'h0950051b03650f520872f1dc07c7fd66f2ca;
mem[944] = 144'h0c8bfa9f08ea0f04ff60fe56f4acfe58fbfb;
mem[945] = 144'hf218f19ffb2bf2d00a290fc60a70fcb808e2;
mem[946] = 144'hfa54fa52f3c2fb72fee3f44dfdf6093c0292;
mem[947] = 144'h0744fad9021a0f1bfa7bf7cbffe7f214f856;
mem[948] = 144'hfd1bfbf1089efd0c0058fb1c004a0bedffa0;
mem[949] = 144'hf8cdefadf227088efb7bf03b050d0c57080f;
mem[950] = 144'h0524f2aefe2702f4f116f330f94d04590b73;
mem[951] = 144'hf23efc5b0fb5f0b6fa9a06f708e90fda07c0;
mem[952] = 144'h028107b4fa61f0d9f9f007f0f42b0b9cf013;
mem[953] = 144'h0974faeb0d20fc750941fd830ee50a8803e8;
mem[954] = 144'h06ea0477f831f113f9faf3b80227fe4c0330;
mem[955] = 144'hfd7c0a8defccf982f110fb8602790d45ef45;
mem[956] = 144'h0b37f2e7f28af4bf09a6f7cff68106c9f1dc;
mem[957] = 144'h094ff453f99006f9fe50f741f1810573fccf;
mem[958] = 144'hf0d2ffa5f3daef650c720252f7380a490804;
mem[959] = 144'h0cfb07b909ffff19eeb90831f4fb0a1ef8da;
mem[960] = 144'hff75f38d029b0f1f0a33031dfe040c19feb8;
mem[961] = 144'h03d80f1ffba6fbdf006907670d640dbbf553;
mem[962] = 144'hf786fb7ef540f9970ef9f973fe540d3a0bfa;
mem[963] = 144'h0948f881f49609d3fc55f8dd0e04f3cf063f;
mem[964] = 144'hf9e3f59c0958f5860681f4e203d9f733089c;
mem[965] = 144'h08580d6f038af2ccf6e3f7c50c15f39b0d2c;
mem[966] = 144'h06f1fbbdffd90e050e3feff1053a04000b2a;
mem[967] = 144'h01840c78fb300eecfa2c024701caf806089f;
mem[968] = 144'hf1d20728f587f73ef8adf2e2fdf4094bf86c;
mem[969] = 144'h0535f5bcf0db0215f4d0f745f421fd1c08e3;
mem[970] = 144'hf50dfa530e890a31f8b70206ff1cf534fb43;
mem[971] = 144'h048001410eb40171f023fc7ef09e0b7f0c28;
mem[972] = 144'hfa44034c0aedf6d20cf9097b016dff74f371;
mem[973] = 144'hf0f6ff56fe1df911fd29090cf67afb14fcfb;
mem[974] = 144'h0f35f56405f3ff9af16bf99704430193f11a;
mem[975] = 144'hf858f6510449fd82f9660dd6f356fa23fb55;
mem[976] = 144'hfcb4077e04b7f7a3f3db011c0867f605f47b;
mem[977] = 144'hf4e1f23ef9e1f45afec3f372f1b60293f147;
mem[978] = 144'h08cef2d0f9790780fc7901e4f647f74d087e;
mem[979] = 144'h07c6033f000a0e250910f4c001330ebd0baa;
mem[980] = 144'hf3e40b8b0abc05d00f1ef1eb00ccf61208ed;
mem[981] = 144'hf2400a530864098bf0710434fca0f85805d3;
mem[982] = 144'hf4de05b803e20a2e00070a9eff440d77f6dc;
mem[983] = 144'hfc1a00d40021fcc10e0604050175fc5808ce;
mem[984] = 144'hfd7700f3fb17fd3c0415f9ca070509510152;
mem[985] = 144'h0b29f9fe043bfe5d035f0d45f472fd0ff2f1;
mem[986] = 144'h0a53f33af0ac0fc00904fd240e930761ff2a;
mem[987] = 144'hfe5707760bc605aef7e2fe3d0b7108f5fc9f;
mem[988] = 144'hf32bf5160723f6db079b0dda087904360070;
mem[989] = 144'hf9c2f323fb3e0090f405047dfb59f9bdf274;
mem[990] = 144'hf99af03ef099f96bfce6f66b04b401b0f57d;
mem[991] = 144'h0f40fc040bda077cfdb70ec0061ef8d6f21b;
mem[992] = 144'hfed6f7a2066bf74af2d1f5cbf61bf73ef507;
mem[993] = 144'h0863f365fdbc00a508e1f9d905ed0b9df9a2;
mem[994] = 144'h05f405abf1dbf6e5ee5af41bfd84ef51f151;
mem[995] = 144'hf80a0678f84a0380f48905adffa007ecf8e1;
mem[996] = 144'h0ae6096ffdc407c3f01cfdcbf3bd0852f281;
mem[997] = 144'h0eedf8240bb9fb39f2ecf2150ac80f990315;
mem[998] = 144'h064802440a8bfe11fe4c08c1fe6bfe5d01c8;
mem[999] = 144'h0f08fd19f18e031807aaf51cf4fbf872f4c8;
mem[1000] = 144'h0b4bf8acf1d50788045f090f002cf9bcf823;
mem[1001] = 144'h08c70bb2fc710afffce6fc00f34b0834efcc;
mem[1002] = 144'hff020c5704360da2f8bdf1030348ffb70960;
mem[1003] = 144'hfd470aa103260eadf2e5f5c80ceafd810ab0;
mem[1004] = 144'hf6adf5f9fcd1fb4ffdf70091016f0b60fe31;
mem[1005] = 144'hf289f59bff95fd36fee606ef057e079ff61c;
mem[1006] = 144'hffd3ef4df536f591f9eafa6ef7ebfebb073c;
mem[1007] = 144'h070303ab0c4ffa9d012efdff0b1cf775f92d;
mem[1008] = 144'hf67901baf4d000760f010765f34df0d607cf;
mem[1009] = 144'hf872faeb0def0254f93608ae0100fe7bfbc1;
mem[1010] = 144'h036008edf4630a320db30a360ebcf8b4fe9c;
mem[1011] = 144'h0b8503680f5cfa39fc510232095af7e60140;
mem[1012] = 144'hf4810b6b0d38f563f5870792fca20a7cf86a;
mem[1013] = 144'heff903cdfc1c01a6023e04240630f9960be4;
mem[1014] = 144'h0c2907daf432f825f7b20772fc9300e4f038;
mem[1015] = 144'hfc86f88c0e17f621f461f785fc230eacf5bf;
mem[1016] = 144'h08860f65fc6b0878fd070c010eccf9f804c1;
mem[1017] = 144'h0074f36af763f043f81f03daf6effec8f513;
mem[1018] = 144'h03fcf7240ba904a4f09c06a0f88b0b9df17a;
mem[1019] = 144'h0c06efd101a1f31c07e9faabef050e06fb7b;
mem[1020] = 144'hf9c50d28fcfafbc8f87400740d1708daf7ee;
mem[1021] = 144'hf897f85a0e420928f80d063c0258f053031f;
mem[1022] = 144'hf6afff64016008e8f0100c81f34602e6f4a6;
mem[1023] = 144'h07050930fa94fa86f8d9f66ff19c0d360543;
mem[1024] = 144'h002ffde3f50cf7e3f19afc16f6a7fad106b4;
mem[1025] = 144'hff9d040c0967f54502a7056cffa40e210336;
mem[1026] = 144'h0d5dfb6808fa09f8f3ca06f3fb2df59d0464;
mem[1027] = 144'hf1f30e87fb6af1a90611fe0106030ee4f9da;
mem[1028] = 144'h0fe50047fd01f0d2f047015cfc7df7be09d4;
mem[1029] = 144'h05c901f6f51cf55d0f880c83f771fc010566;
mem[1030] = 144'hfe47f02d0d7bfa3df5f2011af4f105a40467;
mem[1031] = 144'h044609cdf4ba06fd0b1e0994fdc307bbfbb8;
mem[1032] = 144'hfaf9f2050eabf0620d34f869f3090e1ef598;
mem[1033] = 144'hff400ca40e290b67f53a0c8def3df550f358;
mem[1034] = 144'hf49a0552007bf37e026b03b6097afa7e0284;
mem[1035] = 144'hfa93f0d9febe0127f66ff40e0e7f05bbf4c5;
mem[1036] = 144'h02e40c48fe87efe1f968f05007cdf9e2080b;
mem[1037] = 144'h0778fead022dfcdd088f07c107ebfa30061a;
mem[1038] = 144'h05e90a31ff94fc59f186fd4b00fff6690e5b;
mem[1039] = 144'h0789f9fa08f40406fe07ef480e1b03cef1cd;
mem[1040] = 144'hf48cfd33fd9b0bb109c8efa005bb018f0547;
mem[1041] = 144'hfdf7ffd7fa8a0703060cf4a40e65f80d0431;
mem[1042] = 144'hfc48f0bc09d309acf3b8f1e6fa9f0a2f05e9;
mem[1043] = 144'h03d306130625fe67f11b08b2f5e5ffb6fd2d;
mem[1044] = 144'h017703ae05f30c1e07390e7b056d0e490c69;
mem[1045] = 144'hf19202f70bb2f57b0d0afa6a0739015905ec;
mem[1046] = 144'hef9cfd2e01a3febc01fbf2c70c910b9d0b23;
mem[1047] = 144'hf17df07efe66f429fe46f4b60a92f21201b2;
mem[1048] = 144'h0c7cfdb109fff7a50265f7de0b81f8a2062a;
mem[1049] = 144'hf6920a17f8bffd54f4b9fada03fd06e9efe5;
mem[1050] = 144'hf76904a20a6703f804680968018af876faf8;
mem[1051] = 144'h075bf46f09eff451f72d03640019027cfa69;
mem[1052] = 144'h01b5f5db0066f9c600e909be07a3f639f315;
mem[1053] = 144'h0b94095f0f5df3bcfe010752fa3e05120b02;
mem[1054] = 144'h06b70f030efd0e37056bf617089608010411;
mem[1055] = 144'h0bb4f5240a49022b0c5df06502c505b308b8;
mem[1056] = 144'hf818f97604720ccb09590e54faa5fea3fef5;
mem[1057] = 144'h0299ff59f0b80f95f60efed907c0f0cffc49;
mem[1058] = 144'h0c8f0b13fedb0a86fce5fdae0e50fd52f9ad;
mem[1059] = 144'hfdf7f2d304160142f722f10c0866fcdc0d98;
mem[1060] = 144'h0179fdb90ae704ec0db50b1d04fbf27e0ea8;
mem[1061] = 144'hff61f7b5f3b8f7c6057bfb34f895f33ff3bf;
mem[1062] = 144'hf4f4f00afa2d091cf9f8058dfbb601f50768;
mem[1063] = 144'h06dffe7c0cb7fdf70d8cf593f2f4f4bb03d2;
mem[1064] = 144'h0518f4f50157f4f8f2aafca7ff67f9bdff85;
mem[1065] = 144'h03d2fac60a18f60b0bf30251fa38fd4ef088;
mem[1066] = 144'h0eed0baffd17f767f1f408a0f7a30632f8dd;
mem[1067] = 144'h04b3f598f4060a67effefb67015af70defa8;
mem[1068] = 144'hff6dfe5af44f0f15f1ff0efbf657029ff05d;
mem[1069] = 144'hf2110f2800180fcbf8ee052907ac0be10d5c;
mem[1070] = 144'h0138fb20f730f729fc50f2820c38f89b0dd8;
mem[1071] = 144'hfe22f2fa0d33f0d301f70eb40acb0686f183;
mem[1072] = 144'h095ff848f218f3e1045ffc570019fa0ef975;
mem[1073] = 144'hffb9fd33f78e097afd660c36ff4508a4f326;
mem[1074] = 144'hf75407cb015e06a9f2350d1605ef0fa9fd3c;
mem[1075] = 144'hf70bffecf6960e470b5d028c0595f8d10543;
mem[1076] = 144'h0c27f4fb04f0fe330ef000e3fd4e024c0f04;
mem[1077] = 144'h00ce0f66044702d10a0608f403d60927f02b;
mem[1078] = 144'h0515f6fe09370f7dff5af104072d0e8ef004;
mem[1079] = 144'hfd6efba9f73f0da9fcc60d05f777fda2f836;
mem[1080] = 144'h066ff23b0505f831f2c009d1fd33f39403e2;
mem[1081] = 144'h0a6a03a6fdf0f3c2f20905a0f2e3ff26fea4;
mem[1082] = 144'h0ed804530668f34707c7ef90f8f7f70dfdc8;
mem[1083] = 144'h01340873f344f65901eaf1f005bffb44082a;
mem[1084] = 144'hfcc7ff8b06f40b590263fc3304ccf466fb1c;
mem[1085] = 144'h00620181054402aaf3100d47f360043401c1;
mem[1086] = 144'hfd550c46092cefc3fa87fc45f9ee08080d2c;
mem[1087] = 144'hf10c03090594f8c40251042b02c5f74ffa23;
mem[1088] = 144'h086afb66f630f423fc7df4edf5940572f403;
mem[1089] = 144'h01b7f77d043ef4100c5afa81fc3af26a09ec;
mem[1090] = 144'hffd2f9630aa3f68702e5f395f37ff4130d9a;
mem[1091] = 144'hfb61f57801acf9e8f13c02210260f4fcf726;
mem[1092] = 144'hf53ff92bf131081b100a0b56f97707000468;
mem[1093] = 144'h074ffec2f847f895ffec0eeafa690a92f7f4;
mem[1094] = 144'h07d1f06ffcbef43f050ef5f5f49bfc27eeb3;
mem[1095] = 144'h063b03800b58f9860157f9920982f73906ba;
mem[1096] = 144'h02660abafb51f84f0dc9102ff7c5f71a055c;
mem[1097] = 144'hf3c3fc940d6903b0ffe0023c0f1cfcd603e9;
mem[1098] = 144'h067a0862f98bff13f61bf56808190cbdf3fa;
mem[1099] = 144'h05cb0a91f354f1510795f1b0f15afe28ef34;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule