/*
Copyright 2019, Grant Yu

This program is free software: you can redistribute it and/or modify
it under the terms of the GNU General Public License as published by
the Free Software Foundation, either version 3 of the License, or
(at your option) any later version.

This program is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of
MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
GNU General Public License for more details.

You should have received a copy of the GNU General Public License
along with this program.  If not, see <https://www.gnu.org/licenses/>.
*/

`timescale 1ns/1ns

module wt_fc1_mem3 #(parameter ADDR_WIDTH = 10, DATA_WIDTH = 144, DEPTH = 1024) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h08dff4cb0d5cff3c099af13dfd4e05cb0644;
mem[1] = 144'h0c54fc0900470929fb330eb4f799fe7b0e59;
mem[2] = 144'hf97202d5f56a08c80079f933f7f4060903c6;
mem[3] = 144'h0878f9610d4604c90115026f07c9fc4a0f99;
mem[4] = 144'hfb05098a0ddbfb270bc6f2defe51f8b201e0;
mem[5] = 144'hf1d1fbddf24b0c07fb67f2590494f98ef951;
mem[6] = 144'hf380087af6b8f4cff3da02ccf7560a44f76e;
mem[7] = 144'h0ae80a87f938f60608d3f87d0b16f57cfb24;
mem[8] = 144'h02920bcaf774029402a704ba073ffe29f189;
mem[9] = 144'hfdd5fed10c1df35e0eddfcdefda7f66ff18b;
mem[10] = 144'hf7e6f14200100cfcfb87effbf86ff52c088a;
mem[11] = 144'h03d8f912f11308580bc6f10001ebf27efb11;
mem[12] = 144'hfe5df7660a9b0b330e6e02a3048cfa2d0f4a;
mem[13] = 144'hf8a0038903a9f0f5035ff24bf3fdf2f0f426;
mem[14] = 144'hf7c606590375010c0725f4f1fbc1f071f121;
mem[15] = 144'hf6200bfcfa740e3f06510340f84d0f7ff9a0;
mem[16] = 144'hfda7faadfdbf0fd6f995002607ac04d3f30c;
mem[17] = 144'h06240877fa8a033e0c16f8a304e50386f054;
mem[18] = 144'h0106f533f8c6004902790bc1f83af7dff24a;
mem[19] = 144'hfe810e41058101a6fa4cfa1b0b160c94fa11;
mem[20] = 144'h0f96f66d05e5febef1bafbc90ba60a22fa2e;
mem[21] = 144'h00450f99f244f0dbf11fff3df632fd9b00b3;
mem[22] = 144'hf87100010e39f9c6f3e00b54f46efe040c43;
mem[23] = 144'hfc5efc6ffc22043103720ef1fc83f71dfea6;
mem[24] = 144'h00c4087900aefdee068b03b7f105fa9407f5;
mem[25] = 144'hf4a20e64f38f0f1e0d5d0e5bfa2a0281f253;
mem[26] = 144'h07f40f370409083ef957007ef4160ab404f6;
mem[27] = 144'h00ebff96f061f76af65008c6f591fd08f5e3;
mem[28] = 144'hf18df3270ed9faaff788f4790ed50607f66c;
mem[29] = 144'h01920001f1d00b14ff05f0a0f3930193f853;
mem[30] = 144'h05380eb1ff260948f516f53d0c14f85c0de6;
mem[31] = 144'hfeebfc9cfd470886f23cfe70ff25fc8a03f3;
mem[32] = 144'hf7f40183f28cffaf089a0c560c8bf790f7dd;
mem[33] = 144'h0c7f0cabefea0e4defb00d8bfb10012cf543;
mem[34] = 144'h002cf5a2f028f0c9efc20b75f6b4f883f607;
mem[35] = 144'hf6660736fce50026f70705fef3cffda8f038;
mem[36] = 144'hf95304eb04cefbd3edd9fa8d047301a50e75;
mem[37] = 144'hfe9500feefd6027bf63c06550683fb50030c;
mem[38] = 144'h06eafa0500ff071cfa2ef2c508e6f14ff0cb;
mem[39] = 144'hfdbff909faa0ecc7fd2df1f0fd6405dff111;
mem[40] = 144'hfb97fc1bf95e03d3fac5f2fcfed3f1befec5;
mem[41] = 144'hff5bf9e4069606e8ed4a0a53febc050d07c5;
mem[42] = 144'hfa67fc88ffb8f24c0a13f70501ba011a078d;
mem[43] = 144'hfc8b0b9bf63a0b1a02320d61fe19f7b60cc3;
mem[44] = 144'hf0f5fc460cebf164fc4809d50cd5fef8fe3d;
mem[45] = 144'h01a700b600e6fe6a03ae04150cfdfaa30cf0;
mem[46] = 144'hf944063806420e640dd0f4ebf27b0eb20800;
mem[47] = 144'h04a9f707ef2d09baff2af85ef53e0abcf6b9;
mem[48] = 144'hf9c301600249001c0194fc29f0c8ff420de5;
mem[49] = 144'hfc1205320261043105de0bd7fe43000b0806;
mem[50] = 144'hffee07eafcb80f32fb28019b0294f439fabc;
mem[51] = 144'h0bc208f8f9aafc51ef9af10efc960280fa84;
mem[52] = 144'h0a4b0344f93e0dd0f37af71af965fad1ee45;
mem[53] = 144'hf794fbf1017ef6a0099ff30df0f402d4ee4a;
mem[54] = 144'h02b709d40a9e02cdfbab00a708eff671070a;
mem[55] = 144'hfad305b4f4520affeb72f70a0ae3f067f757;
mem[56] = 144'hf0ff00bef7d10382fdf60d72ffbe0b08f66b;
mem[57] = 144'h0e9d031ef467013c01e30c3c038fef1f09ab;
mem[58] = 144'h06e1fcf1fa8b0d4ef587efc90ef005cafed5;
mem[59] = 144'h0512f73bfb6bff0ffc870430ff6407be0249;
mem[60] = 144'h0730015902b00857f8d90549073e0c62f09b;
mem[61] = 144'hf05dfef9012cf655f40d0d97f1d2f87901e2;
mem[62] = 144'hfbe3f4bf05a1f64800a00c930a70f4ec02ae;
mem[63] = 144'hff920507f43f0a32f04af046f3e6f457f1ed;
mem[64] = 144'hfa70f4fe0a9308940122f8b4f4560de0ff51;
mem[65] = 144'h09730e9ef5290c1efa8df534fbc9f8fc0a8e;
mem[66] = 144'h0c620e38f0d9f7ae00bbfe830ab9fb03f9f4;
mem[67] = 144'h0274f2390dc400ddf422f0de0743f2980973;
mem[68] = 144'hee74f1a3093e0d5afd6806590277efadf76d;
mem[69] = 144'hf8f9f4d0f7ea0564fcc6f7fdedf105ef0736;
mem[70] = 144'hfa7006db0e510241f716f85b04a80b6cf8db;
mem[71] = 144'hefb3088bfb5608d3fe0ef43e06d7f4ce06df;
mem[72] = 144'hfd8fefbdff76f1af0932002af08700590799;
mem[73] = 144'hf1a10701fa89f5d20c49f825f1d6f31c00fa;
mem[74] = 144'h079806f4ef7a069b08ebfc13f17506c9006d;
mem[75] = 144'hf8ea0695f4960493fd1803bcfcd50f55f73e;
mem[76] = 144'h0373fc980c0900170dd7fbd0f06bf571fb74;
mem[77] = 144'h0b7d00b3f085eff9fcf70965022efaa4f0a6;
mem[78] = 144'hf610fe2d0558fc1ef9bff46afd110bff0485;
mem[79] = 144'hfadbfb14fe240e73ffa90b48f661fd4d0d36;
mem[80] = 144'h0937f3befb1bfc6a0760f77cfd92f7b70c3d;
mem[81] = 144'h096ef3e6f62bf3edf9ac0722fa8d0c0b0361;
mem[82] = 144'h075d050e0b590cd5f2f10b320b480823fd72;
mem[83] = 144'h069df56707a3f8970dd8f532f5f30a1e0a07;
mem[84] = 144'hf796085bffcafe85fff304aa02400f2bfe9d;
mem[85] = 144'h06fc0d8a003af1d8ff500e250eb60269f5fa;
mem[86] = 144'hfaa7f0a70f7a0d11f0cf0d84fcfa01c1034d;
mem[87] = 144'hf3aef6d9f46dff8df2c00191fa83070a06a6;
mem[88] = 144'hf29df4b802e3fbcdf27702ee0ee00e94f98f;
mem[89] = 144'h02a6efc40c90052c09d3fe640d8afdaf025c;
mem[90] = 144'h0fc4f7db0ac905a209f6f2a108180161fb28;
mem[91] = 144'hf189f9c1f52ef7d1f5e702250a71f873f04b;
mem[92] = 144'h0209fcd0072701b1fa16093603a1f339f9bc;
mem[93] = 144'hf339f1600378f2f6fb04f76f092e017cf7b4;
mem[94] = 144'h0f6902be07950b1e0c71f6b20dc0fbdef5ea;
mem[95] = 144'h06af0838f29b088307ccfcce0da0f93df899;
mem[96] = 144'hf117fcbb08f2fe8108c1f66a0872f6b008eb;
mem[97] = 144'hfb1b0474f4a30a0804bcf58ef8830dda007d;
mem[98] = 144'h0cbd0167f68efe59f8b6fb21049a0c74f2ce;
mem[99] = 144'h096701aef948f4befa28f54d040ffd6bf9da;
mem[100] = 144'hfb41fdbaf823fbc5f7e9f3250640eec7face;
mem[101] = 144'h08d3f3befba40e0ff5d6fb9605070390f53e;
mem[102] = 144'hfebc0928fb7b000cfb90fcb2fb02f5aa087b;
mem[103] = 144'hf44909180426fa4bf674035f00dbf9c1ff67;
mem[104] = 144'hf606f51af60def3107c0fcbaf073f825090d;
mem[105] = 144'h0eacf9c703c3eebf06cbf0030e6d000af950;
mem[106] = 144'hf9e5f7b7fee0013906cd0052f99d02100d98;
mem[107] = 144'hf3c80659f1e1068d061103820280fce70496;
mem[108] = 144'h0d9507defd33033afe5008e7fd21ff7303a6;
mem[109] = 144'hfae3f8ef027cf2490c92fa1ff1350774072c;
mem[110] = 144'hf18af8d9f5e8042708d2011ff94ef8bcf622;
mem[111] = 144'hfc35fa4af1d5fc070bca00a9f45d0bc7f35a;
mem[112] = 144'h07000a5a06a3f43c0cb6fc1800b1f8b1f08f;
mem[113] = 144'h0d00fbd400150f480d62f327083b09890e02;
mem[114] = 144'h097d031f0b87f1f402d6f7940f8506bb01ea;
mem[115] = 144'h0145ee12f9f70b82fec8f33ef7930b540c0c;
mem[116] = 144'h096b01cd07bdfa45f4a90dc10351f400f493;
mem[117] = 144'h00bcfa7e0267fbde0c2404000cff004c0744;
mem[118] = 144'hfa0f0715003f08bd00e4efd3f294f19d0dd9;
mem[119] = 144'hff87febdf20f072001f304acf8d1088eed67;
mem[120] = 144'hec4cf084fdedf4b4046709190468f6c10eec;
mem[121] = 144'h0c120ce3f43105d2fba001fe070e0e18f000;
mem[122] = 144'hfec003810e2a0f7a0dea0094f16dfc50fe68;
mem[123] = 144'h03e7f155fb3103a60632f209fdcaf6ac06f4;
mem[124] = 144'hf4fb0c82f1fef6d4fdb4003700560090fb18;
mem[125] = 144'hf63c06f8f2fd046a007fff80f4a702d7ff89;
mem[126] = 144'hf8f3f43df972fa5e03810844f9ea05ac0077;
mem[127] = 144'hf718fb7ef8ccf3ac0aa0f65bfeeffa83f896;
mem[128] = 144'h0be8f5ea02e70845f46b0307082308d308a8;
mem[129] = 144'hf93201f5f082f7660c94fa0cf7b00efc07b0;
mem[130] = 144'hfe55f781f1cbf32cf025f19f0f53f7e3055d;
mem[131] = 144'hfc8af8960219f5fcfbc4f89e05d908930412;
mem[132] = 144'hf4fff95f0900ff9b077a0e16ff680558fc4a;
mem[133] = 144'hf96a00f1041e0a7df52f08960c4cf4f7f887;
mem[134] = 144'h0739061204c409b5f941f76df2bcf5fbf818;
mem[135] = 144'hfa3903220cc2f483ffaff761f2c70318f89e;
mem[136] = 144'h081e014bf35b0883f3c20e98fd0d00290bde;
mem[137] = 144'hf8a307330f4b0e0d06c2f838fb3d0fd0fa45;
mem[138] = 144'hf6950c4b02b9f3f708610c94ff85fb1b018c;
mem[139] = 144'hfb080e8f0f7b0e110c71f5cef80b0931f9f0;
mem[140] = 144'hf03dfb99fc1b025a0708f26ff8f7017505e2;
mem[141] = 144'h056bfc7606dd0176f326feaf031e09c6076b;
mem[142] = 144'h0e4d0673fa2607070885fc520f250ca60266;
mem[143] = 144'h090af4e1f429f8c7054301ae009efdfdf0a2;
mem[144] = 144'hf9180000fc0702150967f88ff567fa9105ee;
mem[145] = 144'hf516f63afee50d350fe7fb200ea700a7065e;
mem[146] = 144'hf7820a3bf727fbc7f0f5f44d05d8fe71f3b0;
mem[147] = 144'h0306045d06b7fdcf04abf531f93af65af1d7;
mem[148] = 144'hf699f6930e3e0b2bfc95087b019403290912;
mem[149] = 144'h0534f2a8fa3af891f88002eb0e03f09909e8;
mem[150] = 144'hff54ffbcf48104bcf033075cf5860e8afd05;
mem[151] = 144'hef9dfd6cf108f40a0da1fc55f61bffd90724;
mem[152] = 144'hfcc50e05fb4bf43a080f0e56fb39fe23fa48;
mem[153] = 144'h04410b9e0145001ff1bcf9710675f8170e1c;
mem[154] = 144'h08d6f77ef7fe0c7a04bdfdc10f47f5d7eff5;
mem[155] = 144'h07befee40759f560f4e2fae4fd5600d90283;
mem[156] = 144'h06befb42f47f07b80a630cd5fdd103d1f98a;
mem[157] = 144'hf033f948f73e00d4019803790588fd58f108;
mem[158] = 144'h03b1f3ca0b4bf4dcfcb1038df5d3f05305ca;
mem[159] = 144'hf76f0b44ffad06fffcbb072200a0fb87009f;
mem[160] = 144'h0504f40afc9a04c1f60f03eb0586034c0bc3;
mem[161] = 144'hfe85fc99f17905a4f255fcc40d88f39807d4;
mem[162] = 144'hf224093bf172006efc0d028009220dccfa19;
mem[163] = 144'h057bf653fd16fb9efee6f1170e1bf47505b2;
mem[164] = 144'hf4f00c870f1af22e007a03da0978fd4908fc;
mem[165] = 144'hfcc3028b0e82f070f017f597f314f4340fca;
mem[166] = 144'hf1ccf639f2cf032bf8e40ca30d5bfc1ef0cc;
mem[167] = 144'h02ea0513088e0c27f0a6f41ff1f6f20207d3;
mem[168] = 144'hfccaf93f052afdfbfa6eff99f82002a104ac;
mem[169] = 144'hf432f2bdfdc904b202b8f2a708d5f96c0984;
mem[170] = 144'hfc39fab2f22bf0cd0293017803450909f9c5;
mem[171] = 144'hf96df733076d0557f87ff3cef171f9ea0ffb;
mem[172] = 144'h04a40836fb3400dcff8b0703005cf846f368;
mem[173] = 144'hf257ff2007e5f6d5fa5c05a10723fc20fcd9;
mem[174] = 144'hfcbaf8d90ba30cc1055cf1b1f479fe62fae2;
mem[175] = 144'h0f73fb9ef070f372fc220dc8fd0cf04ff7f3;
mem[176] = 144'hf76b0ba9fdb40989f0ec09b803c9f5e20293;
mem[177] = 144'hf7c1facdfe1a0733f424f915f8c404be0bf0;
mem[178] = 144'hf91702d90808fc29f54b0cf0fb2803b30f62;
mem[179] = 144'hf042059c03790c310c7ff21cf775f362fb6b;
mem[180] = 144'h01ca0334032900d606ab0e41fdf903b604db;
mem[181] = 144'h011ef302fa710234fdbaf0610c6cf89dfc62;
mem[182] = 144'h0f3c0519f7d2f98703e7074208a0073ffeee;
mem[183] = 144'h00c9049fef64fe810cc2efa90ead0daa04f9;
mem[184] = 144'h09b9ff40febffb23055008abf9520aadf7cb;
mem[185] = 144'h070ffa1b05220172037ff3ff09fef95efe75;
mem[186] = 144'hf77e02f4f291fe1ef92f02d80a2d04c70186;
mem[187] = 144'hf683ffc8098a01f7fd620b92f690050bf187;
mem[188] = 144'hf50ef24004aff112f71cf54df6acffc60bde;
mem[189] = 144'hf2c7fd42fd74023309cbf666fbe90106fb02;
mem[190] = 144'hf6040fa8fdc60abcf85afdeaf631f599fa29;
mem[191] = 144'h0598f947fa6df2aa02a90b4ef4f7f4c80f50;
mem[192] = 144'h038c0885fd86f70df413f345f033f2ca0404;
mem[193] = 144'hefdefb3af51c05f10f69fa09f6f8f5f20eca;
mem[194] = 144'hfdbefdf50656f00df9c9088508f9f8430c59;
mem[195] = 144'h0622f1940e760993f829ef3d0518f59ef487;
mem[196] = 144'hf3a5f4deefb2fa790f99f332f6fceee8faf6;
mem[197] = 144'h03ac01a80410f0c0fb26f4ceffe1069a0baa;
mem[198] = 144'hf1e6f4f6f4300ed7f778f84b0a80f38e03f8;
mem[199] = 144'h00050a92ee0af871f432fd77fbc7fdce06cf;
mem[200] = 144'hef78f7ebf437f83afad2f905f86cfc020bdb;
mem[201] = 144'hfdb1f51afd7d08b6f911f2d200b2023a0c1f;
mem[202] = 144'hfdf7f23a0516f062f12a0d9afd56fee5f856;
mem[203] = 144'hf912fca80a1002a00e5ffccdf72af33cf8e9;
mem[204] = 144'hf17208a3fbd3f739fdf2ef64084ff1320cd1;
mem[205] = 144'h0af3fa2503e50f5906a1ffbb0ad10b70f96f;
mem[206] = 144'hf3e9f3830f3501090322f850f3ddf92b0d90;
mem[207] = 144'h009d0e2904a9f435f92e099d0440fc0af651;
mem[208] = 144'heffc01eef6e70b64f3f7070407a3f9b7f379;
mem[209] = 144'h026bfb9f01bc097cf2b405b5f72b0b180f42;
mem[210] = 144'hfe1301960d6606f6f89e0685f17b0431f0ba;
mem[211] = 144'heed0fc8608b8eed403f3018ef301f60df075;
mem[212] = 144'h0127ff71f45bf9c9f07704fc0468fac8f89d;
mem[213] = 144'h0333fe00ee1c01fc0e33ff6a07eaf9affe6a;
mem[214] = 144'hfb92fb3805dc0c43f3e707a00eb60224040d;
mem[215] = 144'hfb7bffdbf707fbf908a5f7cc054b06330039;
mem[216] = 144'hfbfbf99ef080fcd6efed06d8f6240878fd10;
mem[217] = 144'h0052fdc2067df70ffdb9f79ff460f6adf4c5;
mem[218] = 144'hf024064307f805e3f43ef4640a7102d0034a;
mem[219] = 144'h008d075b0489f231061d09d5f097f5f8fba0;
mem[220] = 144'hfd910763076bf959ff7df244f405f52e098a;
mem[221] = 144'hf134f53efab3f78008130da3f3bfef3d0712;
mem[222] = 144'h0696facc0884f8fffca100010030fb7afb81;
mem[223] = 144'hefc3fbf2ffc5fb2a046d07430ecc0a65f71f;
mem[224] = 144'h0dfcfc65ffe50cf3f41b04bd0fb9f75ef6d0;
mem[225] = 144'h0490f3720a1a00f205c80d43f7080e040d58;
mem[226] = 144'h0ec0fb490d15fb0af9d3fd83fb4a06410ba0;
mem[227] = 144'hf5aef309fb1702b1002bf730fd30f66e09c0;
mem[228] = 144'h0a5cf200f6fd0752fe720659fb1df795efe8;
mem[229] = 144'h033f093e09960350f7e7f876065af243f0a4;
mem[230] = 144'h076af478f05004c10838f6550799f75b0004;
mem[231] = 144'h0c15f4e6f8b208a4ffadf01203d5fd77032d;
mem[232] = 144'hf40502ee00600e26017c01fcf89df86fff9f;
mem[233] = 144'hf37bf61b059fee42fb0409e9f694fe12f469;
mem[234] = 144'h0a58fc10f63e04d4feabf0b7f479f0050f95;
mem[235] = 144'hff6902a9f339f873f40ffbc1f8adf4b1fb66;
mem[236] = 144'hef92f676f26f02f7f34105e904f704aa0d33;
mem[237] = 144'hf037f54b04540ad6f8b3099306f4fa240bca;
mem[238] = 144'h07390550fb33005d078a0fa7f4e40849f82d;
mem[239] = 144'hf3f20bfc0aa0fc36ef8c0ad6099900f7f8ba;
mem[240] = 144'h036dff7bf13ef9570de5ff1df4020d17f127;
mem[241] = 144'h04d7ffa8f2b008260db6f2abf77ef316f8f0;
mem[242] = 144'h0da90fdd09c604f102a60e9efb6cfceaf7d6;
mem[243] = 144'h068eff96f83cfcc2f11bfe4403dbfd440bcf;
mem[244] = 144'h047cf095f6560a8cfef50535fb89085e0ac0;
mem[245] = 144'hf60101b2fa29084bf5cef5950b9a068dfc66;
mem[246] = 144'h05abf156039ef5710a9400d8f112086efc79;
mem[247] = 144'hf890f331fb9602d2fcb70692fceb0473038b;
mem[248] = 144'hf99806e5fbae05ff08e6022b0770f44ef2e7;
mem[249] = 144'hf9cef3f60379fc18ee9503930087fabff31d;
mem[250] = 144'h0be10d3bfd7c014ff559f50701a109e60c12;
mem[251] = 144'hf167fd7400a9034a0ce00b1afe80f80ffc35;
mem[252] = 144'h089bffdf0d86f2baf6130c610a00fbbc0e85;
mem[253] = 144'h0317f2720016f58ef8b2f66b00eefc77fcbf;
mem[254] = 144'h0eec050dfae90519fae2f81ff520ff1d06ae;
mem[255] = 144'h007cfc50faab089bf3f8fa240b9c096a08ae;
mem[256] = 144'hfc3d0c5202020739f8bd0dd1fb7f0decfe33;
mem[257] = 144'h057709dbf740001cf489f8ebfd6df951f1c9;
mem[258] = 144'h031dfbad0ffdf56a01360829f424f631fde0;
mem[259] = 144'hfc2df6d809d9f0f8058ff4f9f1d1f935f005;
mem[260] = 144'h0353f483060806a1fd7f06a4020409d4f1f9;
mem[261] = 144'h0d93f5850c120064f201fec6088303d0ef6d;
mem[262] = 144'hef8105b30ee3f5a004dffa33f016f97201e7;
mem[263] = 144'hf6fcf358f278ef7f057ef667fbb50c54ecec;
mem[264] = 144'hff620fa6013f0f0301ed06c6f6ea072d05a7;
mem[265] = 144'h004a093df0ebf53605d506f303d3efb100b3;
mem[266] = 144'h0e0c03c504b1065cfa420ce60e70023e0bd8;
mem[267] = 144'hfec20e38f8c5fd2ef5def8ccf4f90a3f062f;
mem[268] = 144'h0339f8b6f559f9a6045bf4630b770164f87d;
mem[269] = 144'h0485f5f904c9ffcc0dd6f2c9facafb09faaa;
mem[270] = 144'hfe2a0c1f00aaf84bf66c0962fa3afe9303d9;
mem[271] = 144'h0c80fad7f7b7f31cfa450b17f3fff538fc92;
mem[272] = 144'hf0f60cf5f192fadc0e2af314f61df104fa73;
mem[273] = 144'h0b2ffaf1f7dc0d060c4d03130a6909850a44;
mem[274] = 144'h02ad0eea099f03e0094dfbb50f6ef9d3f455;
mem[275] = 144'hf003f50dffbafdd6f98a09e600520a1ff7fa;
mem[276] = 144'hfd2cf74604c0f50fff960359f0860d7d05e5;
mem[277] = 144'hff3ffdc9f7d6ff22f468036ff70f04450ccd;
mem[278] = 144'h015af21f02bbfa62f715057409d5f94e0269;
mem[279] = 144'hf6820808f1aa0db0f03500cb09a6f2d3f78c;
mem[280] = 144'h0a75f0a10e2ef4460211fb2a0051f1f00369;
mem[281] = 144'h00c2fed802c5fe49fbd2f3f702a9fcbdf8e5;
mem[282] = 144'hfcba004c0e60f751f5d00f850bfa0eac0820;
mem[283] = 144'hfb5bf14a06dd0180f951fbbc0ef5f3ba0765;
mem[284] = 144'hf761014b0f25047b0b76fe05f29cfd120b18;
mem[285] = 144'hf16af0f00a390425fdbf057ef87cfd2cf97e;
mem[286] = 144'h0dcef85d0691027afdaffceffb55f873f926;
mem[287] = 144'hf3f2f33efc3902a9f18cf7de0bad06cc005a;
mem[288] = 144'h0afcffe00be8f8b9046b032606da02fff931;
mem[289] = 144'hf08effb4fb27f3f4f027096c034dfe05f5a4;
mem[290] = 144'hf36af0c9fa55fd96fbe5019efd4d062cf6e6;
mem[291] = 144'hf5a2fc67fe59fc8ef1e5eeebf6d9016bf112;
mem[292] = 144'h032201720c080eea0e17f21c03ccf7a700bc;
mem[293] = 144'hfd4cfc55f1bffa1b0d0a08d6f395003afb30;
mem[294] = 144'hfc7101f8ffec03fc010804eb05590bde07d0;
mem[295] = 144'h086beddd0847f247ef39f61dfe960943f5e8;
mem[296] = 144'hfa430ba70065ef04f40f09f602eb057bff99;
mem[297] = 144'h013f0cc9f62bfefd047e065e04390196ff78;
mem[298] = 144'hfb2305b906c7f4e70a74f7f6f9130e4e05e6;
mem[299] = 144'hf3d8f69af73a0871039e0b79f9dff7fdfcc3;
mem[300] = 144'hfa2c0571ff97f498f1d5f8b603a7f5bf0311;
mem[301] = 144'hf34ef009072df1e0f87105fd0b3702f006ab;
mem[302] = 144'h005908ba08b4fa72f95d077b0d4af55b07a1;
mem[303] = 144'hf8fa09b6fc5cf52f03750a8003dc05aa0017;
mem[304] = 144'h02dd00cb0b82f5720be9f76bf5acf165ffe0;
mem[305] = 144'h04b6f351fcf40b45facb08a1f5d3ff7df100;
mem[306] = 144'hfcb608e1f0cd05aa080df715fd01042b08ca;
mem[307] = 144'hfb2d00eaf3ef0c00fe56ffccfb920b59fa6d;
mem[308] = 144'hfa4df4ecffcd01b2f13500dffd0f0bc2fc63;
mem[309] = 144'hfe150a7cf83bf88b093402e5075af74defbc;
mem[310] = 144'hf94c0dfef4bcf8e70e1301d60d0efa0df394;
mem[311] = 144'hef50ec55fe1e05b6ffbc04b0f7afecb8f73e;
mem[312] = 144'hf60905e4f2020679fd14efb4f71c023403fe;
mem[313] = 144'hf8a409dbf66e0046f141fd40077c029a01f9;
mem[314] = 144'h0be1f26ffb1bf4fa0b3a0e84fb9906360591;
mem[315] = 144'h06ebfdd1f44df6ccf1c3fd4ffdb8078805bd;
mem[316] = 144'hf83df0e9ffa6f70dfedef34cfe26f874ff65;
mem[317] = 144'h05e909b106c80b42f6be0464058907f4f7cb;
mem[318] = 144'h036e0bbb0f08fc5bfe32fabb0aad099206f8;
mem[319] = 144'hf0f4f3bbf75ff55d00e3fb4b0439f78ef1ee;
mem[320] = 144'h09990ccffacd053ffbbcf0f30f86fd96f5c9;
mem[321] = 144'h012c01fcf377f599f70d00790935f0a5087a;
mem[322] = 144'h0e0afe140773f5b804dff82f090bf7fef2ca;
mem[323] = 144'h052cf830f236f5de03f00b9601d20662fafa;
mem[324] = 144'hfb75fa72f7d8fe83ee28f8f40714f14cfc3b;
mem[325] = 144'hf2470572f8650a6b0ad0fba70da3f0f0fe64;
mem[326] = 144'hfea4f28f04b4f8f8f8a904a609e8f34804f6;
mem[327] = 144'h07aef4af0b4808cffc71ed5df53e0a5eeddb;
mem[328] = 144'hfd98ea9bf4a2f4790d81f3990c48f0350eaa;
mem[329] = 144'hfef0f91cfca90461f15808fa0168f4b0fecc;
mem[330] = 144'h0f99f1e2fd160135fbb706e4fef908c0002e;
mem[331] = 144'hf58b0623f816034809f2f12a06b80f920f5f;
mem[332] = 144'hf7910dc10a5c0b51078cf3a9f814076e0b3e;
mem[333] = 144'hf9230a27047208d8029d0d31f693fb71fdc8;
mem[334] = 144'h04c5fe6df004000efac3f008f272095af192;
mem[335] = 144'hf9dff8960f27f9420d110bef091906d507e4;
mem[336] = 144'hff9c02680f1b0123f764026ff07c00a50dd9;
mem[337] = 144'h0592000afcba08730f1ef0a20efc02360133;
mem[338] = 144'hf6d5042dff210c4d01780774fddcf163fccf;
mem[339] = 144'h077505e7f8930ea5081006ae0eaa050005d8;
mem[340] = 144'h080201ef021ffc4c0e76044df83ffa5604d8;
mem[341] = 144'hf290fad20216f5ee0aa0fdef0ba8fae5fd5c;
mem[342] = 144'h0f59016005ff0c07f3560c0b01c700890acf;
mem[343] = 144'h083ef126fd540627fc02f9aef69bf25ff877;
mem[344] = 144'hfe330d4b07b7fa790032fb23f2130d2f08b2;
mem[345] = 144'h093afdaeefa9ee5eeeea03170e7f0744098e;
mem[346] = 144'hf4fcf431f4f8f240f3100d89fac60033fd4f;
mem[347] = 144'h0134fdd8f6dd01800bc90d62049cf46ef940;
mem[348] = 144'hfe030df0f087fb47fd9efed2f158fe010906;
mem[349] = 144'hf71afd0af02bf0fc0947ef99fd62ff7c048c;
mem[350] = 144'hf5110a550a83f06600ccf6e30ab7f755fde6;
mem[351] = 144'hf1def1c706330c68f325fa93091bf4c00101;
mem[352] = 144'hf02408cd0e8d0a88f5fd0af2f1460ae40e15;
mem[353] = 144'h0c50fb5505a1feb00a7e04baf458023efa9b;
mem[354] = 144'hf574fa0cfc90f51e0b3afa180270010102e2;
mem[355] = 144'hf65bfa1d0f30001209c7082af0a20b08fe0c;
mem[356] = 144'h0285f4f5f561f2590caff99ff3c403b1f56b;
mem[357] = 144'h04ebf3f401bbf403f69cef27f4f50ceb0a0b;
mem[358] = 144'h0e65f42c02a40f290763ff86087bf6cbf907;
mem[359] = 144'hfd06f0ee09b30194f93ced9f0028f051f0ab;
mem[360] = 144'hf1e5f5f0f123f7cdff0ff169ff7c0eb603ca;
mem[361] = 144'h00490c91f072f13fff61fcbcf4fff712ffba;
mem[362] = 144'h0d380284fa140dd8fdb2f7a5fc270dee06ee;
mem[363] = 144'hf6df0150013b04b70e50f5f3f8b605330e80;
mem[364] = 144'hf618f34af839f71bff74efc4fae203940952;
mem[365] = 144'h0764f61e0c490a9ffb61fbeff079f09efe81;
mem[366] = 144'h0426f65c0748fe200f3d069cf977fd9b0b6e;
mem[367] = 144'h03c10f79f9bff518f25ef266f840f8140ded;
mem[368] = 144'h0d6405260fa1f88e016c01c309bb03f802ea;
mem[369] = 144'hf8780b7301580364096b0b270b330797027c;
mem[370] = 144'hfb190d7f0b85f321fd9afd8304d0f5a3f649;
mem[371] = 144'hf0a3f114f25a0a2bfd5efb54f80cf40c0c19;
mem[372] = 144'h0e3c01b9f17bf8c308e5f9f80208f4a0fbbe;
mem[373] = 144'h0af700d005c801a20598fd95f448f05dffa7;
mem[374] = 144'h09e6f35603110b210d64f8350b330cc90866;
mem[375] = 144'h0b1503b6f431f391f28805f80509f9d7fc88;
mem[376] = 144'h082b0dc30475fcd7f5fc0887f0dc000d0bff;
mem[377] = 144'h0a29f5b10e6a03b9f43808d90b03ff370ebd;
mem[378] = 144'h0f83ffe0f4b1f4b00d620452f9ae05f2fad1;
mem[379] = 144'h09cefef50477fde0fb280f3f0029f3f3fead;
mem[380] = 144'h0f54fb2e04e009f206b1fed60e7af77af201;
mem[381] = 144'h051ef24700a00b5e0e260df4f656028af5e6;
mem[382] = 144'h0c2c0a250d1ff082f3040c31f2660dfb06d2;
mem[383] = 144'h0f59f13bf5dff102fb83f72904d7fad40676;
mem[384] = 144'hfd1fff07f509f5a3f8290ae00b80f824f006;
mem[385] = 144'hf21afad9fb59fba60ccef217f793f2630b58;
mem[386] = 144'h03d6f725f1d6085d026107f3f10e00b3064c;
mem[387] = 144'h0dbafc80f812f672ffe40e75f93ff3c7f67d;
mem[388] = 144'hf8830411f661fbadf23cf664f75af1830841;
mem[389] = 144'hf3f6f01af40f0580f911f48afe60024ff317;
mem[390] = 144'h0e880959f089ffc9fb9a05aefc3ffd3eff30;
mem[391] = 144'h05530847eebb05be00a0ffff0038ef7df880;
mem[392] = 144'hfcd8faddf55209f1f86efca300edf48af6cd;
mem[393] = 144'hf27005d10b6a0adffab8f671fcdef411078c;
mem[394] = 144'h093ff4f3f57cffccfffe038ef1fb06f5f32d;
mem[395] = 144'h0c200a5601ec08defdddf4d30f20f7acfe5d;
mem[396] = 144'hfa4efaea0df60af704aafd7ffdae043e0397;
mem[397] = 144'hf8f2fd87f9b602ef051d09f90169f6db03a4;
mem[398] = 144'h0de8f014ff40f345f1d40eb2f94306e3f63c;
mem[399] = 144'h0495f6c8fc7d01e401c70bc30b6b0e49f180;
mem[400] = 144'h0725f6dff012fdc9f9c3f66f02100cf10cdc;
mem[401] = 144'hf93afe1a04f8fcdc0897fabdfcd208f6045d;
mem[402] = 144'hfdecfbfbfc4e0c9a0893fb4cfced0be102f9;
mem[403] = 144'hfeb5f8cefab6f584032dfa09f54ffd80f25f;
mem[404] = 144'hec73018108ca0914fbdcf999f03ff175f0a6;
mem[405] = 144'hfcbef1dbfa35faaf075ffd0d0ae60aa107aa;
mem[406] = 144'hf9d00ba307a90baff32209a3f2cdfed8f4d4;
mem[407] = 144'h0159eb510653038ff3950a2b0705f5d6ffcf;
mem[408] = 144'h0209f4b9fefcf5030b6efe81fa59f40cfc5c;
mem[409] = 144'hf69af80c0818f45a089705a1fa45fc6904a5;
mem[410] = 144'h09fff574fad00bbaf43c0299fdcbf6110f9b;
mem[411] = 144'h01f50bea0e92f39008800afaf5570db1f780;
mem[412] = 144'h0adf06f70e14f0c5f6fc0954038dfdeff1d0;
mem[413] = 144'hf62a0613f475ff00f8b10809eff3f8a8fea5;
mem[414] = 144'hf74d059e04950393fab7f08303b2f2f70fa7;
mem[415] = 144'h0615fe8608baf257f489f4f901a8fba10724;
mem[416] = 144'hf3ca02cef7e4ff35f06d03bf0816087705d2;
mem[417] = 144'h079af6a8058607540991f62ff8f2f59cfd47;
mem[418] = 144'hfd48f9dcf489f7eb013cfe470eae03a2feda;
mem[419] = 144'hf193fa0203540b0b05520a2b02f4f84bf674;
mem[420] = 144'hf7d4f79ded63eef6f7a9f924fb7ef0cf0014;
mem[421] = 144'hedef01ce029e04ae0878069bf35000650ae7;
mem[422] = 144'h0ab9f78f04df05cdf3ba0e0afd3af17407df;
mem[423] = 144'hfdd4087af4c4ff840416fe7eead1f9cbf043;
mem[424] = 144'hf0d4fc5cf688f248edb1faf3f302f20c0de4;
mem[425] = 144'h05d503d90a63fb00f235fb9cfa720c5e0b18;
mem[426] = 144'h0187f51f0705f9f1fe8c0b8e0161fd610615;
mem[427] = 144'hfd5ff03f0844fa0e075903f5f3e1f3e108e3;
mem[428] = 144'h0cee09c6025cfebc0b3cff9af9ebfd4bf3e4;
mem[429] = 144'h051beeb4f2f70110eed009160a850d99f9ee;
mem[430] = 144'h03640a53fbdbf5b5fab009abf3ea0dc90411;
mem[431] = 144'hf7f3fb26f6a8f5cefc550c5503140a71f040;
mem[432] = 144'h0a12f5e4fb14092002ccf590009d01fef25b;
mem[433] = 144'hffbe0877f4320e90fa46fdcffdcf00e20176;
mem[434] = 144'hf920f135f176031c0f7ff113030ef8aff7b7;
mem[435] = 144'hfb45f17cf2f70751fd0c075606bf0556037c;
mem[436] = 144'h0b2df0ab0e86f7470f5efec00a2dfc8307f2;
mem[437] = 144'hf2b4ff600b4ffae209260144053306be0b26;
mem[438] = 144'hfbd101f4f0360e690b9e0bcaf6de0eb20eb7;
mem[439] = 144'h0cd7efcef5890d48fe3ef7f60ba7f4c9f270;
mem[440] = 144'h051d0d9104c40a91f5a10596f796fe770508;
mem[441] = 144'hf1a7fbd9fbb50ef7f60f07f804acf7f70b91;
mem[442] = 144'h0553fbfef9f2f1220d86032609ac0fab0095;
mem[443] = 144'h0464f921f1ed0edb0847f9a70cacf2e00ad6;
mem[444] = 144'hf3fdf890085e068b0aa2042200c2fcf1f907;
mem[445] = 144'hf5bc0137fc82f289082ff25200dc0d89066c;
mem[446] = 144'h0f0106ccfd8806d7ffd3f3e50b81fc170bc6;
mem[447] = 144'hff3afe1f0578fea2f688fd21f9910272f87d;
mem[448] = 144'h0cf2f62df771f4240e96f91002ab0caa0fdc;
mem[449] = 144'hfd06f842fdfd0c1e07b9f9a1fa1d0d2bf5b8;
mem[450] = 144'h0cf0035d0655f26ef35107400ddb0b58fd35;
mem[451] = 144'hf751067af00406c3f9b6fc14fffdf5eb024b;
mem[452] = 144'h0dc50655fb4b053d0c3af672f3e10d8f0336;
mem[453] = 144'h04180e9efdf0096c024eeffbfd4e058ff3a2;
mem[454] = 144'hf45def520474f73bfe50fb21f2c4fe79f714;
mem[455] = 144'h0c5406760b4602640aeefa27001b0614f52c;
mem[456] = 144'hf19b0356fb6a04b7f6c0f3a600fb00530223;
mem[457] = 144'h050505e104a2f34cf49df280fdaafc7bf47f;
mem[458] = 144'h0346f98700ebf7c200e800db000afb42f265;
mem[459] = 144'hfa9af1d1033f0b38011df007f5d1f2b0fe7b;
mem[460] = 144'hfc310ba1f8c101330dc309b6fd6b071300ff;
mem[461] = 144'hfee1ef1ef171f92d0cb6099d0e5ff7ddf2e3;
mem[462] = 144'h0a1efc4e09f90e2dfe01fba6fe3af5f7f4ba;
mem[463] = 144'hee5bef77fc10f5cafb87f283fb2600600668;
mem[464] = 144'h08830b6d0829f1a30b31f094f618fbc0fa0c;
mem[465] = 144'hf4dd00750de1038105340ea4f2d80f60f786;
mem[466] = 144'h05d60abf0d3bf887f9a103e20dfcf50908a7;
mem[467] = 144'h00e5f151f927fcd9f9f3ffc1f1acf64800b9;
mem[468] = 144'h07dd07d7f400f11df0400ba3f58a00ea03ca;
mem[469] = 144'h0cff045d0523049ff3f9f7f30858fae0f13d;
mem[470] = 144'hf796f96af45a0d7ef62af1d3f1d6f52ff183;
mem[471] = 144'h036ef1e7f3f2f414ee70023feef7eda3f68c;
mem[472] = 144'h06c10eacfce4f6d606da02f7f15f0998f94a;
mem[473] = 144'h0baff1d50e7804baf613f937ef3103aa0398;
mem[474] = 144'h0a98fdc4f886fc240b200bc6f61afa4a0d07;
mem[475] = 144'h0d7a0f5cf5d10bd608f60e2bf2250953fd6c;
mem[476] = 144'hf637f081fc0d0a88f527f7330515f269f71d;
mem[477] = 144'h05d3f528fae20c77009cf5b5ff6cf42ff5c6;
mem[478] = 144'h08cff054f47d07070c2b07bf082702890636;
mem[479] = 144'hff0d04db04a5f460fe5ffe91ffa80f64f441;
mem[480] = 144'h0836f402f7380414f03f066b0019facd09e5;
mem[481] = 144'hf86e00c4021e0ef7f93ff42805750f11f67d;
mem[482] = 144'hf35402d2fc460b15fc27f404082ff84df121;
mem[483] = 144'h03fff8dd0dfc0718fec5fa9ff485030d0467;
mem[484] = 144'hf5a1099d01760929ff1ef184f2d9f8600277;
mem[485] = 144'hfe310e96f294fadc0cfcf12f02f6f4620394;
mem[486] = 144'h02130cc204ae081ef80202a8ff90f187f35b;
mem[487] = 144'hf3a20cdcf7d9f4a9f5c8029c0e320486f01e;
mem[488] = 144'hf07e09a3f21c046af7a90485f6540afdf03e;
mem[489] = 144'hfb8604ebefddf053018906830464fd0af1b6;
mem[490] = 144'h0cd30c43009d0d0ff84afd98fd550c06fedb;
mem[491] = 144'hf772fa98ffc9f8b50aeb021308d7f4260479;
mem[492] = 144'hf98efe400078f333f17ff8370f1f0bad0985;
mem[493] = 144'h0c26f049fd35f14a0e6bf3d7f12ff478f552;
mem[494] = 144'hfbcff67af7c6f706fad9f3ed04b203f702d8;
mem[495] = 144'h0cfcfae9f1d6f6050f4a07cdf681fc590f14;
mem[496] = 144'hfcf604a8fe59f0ee04490e76f1a103cdfec4;
mem[497] = 144'h05e10bf1027c044afac7f6f2f194f9c0f84e;
mem[498] = 144'hf2abfba1f7c705e3ff20f6e5013e05750371;
mem[499] = 144'hf3c7fd530cf7fd550537f3a705de03970846;
mem[500] = 144'hf12cfc34fd3105220cb9fe540890056507af;
mem[501] = 144'h0eac0c25f1d5f29afd89fb3cfd80f509f319;
mem[502] = 144'hff0102fdfa9d0515067e054ffc2409d209a9;
mem[503] = 144'hf0e9f0680d94f7b10203f2df0c1d068cf792;
mem[504] = 144'hf92dff6afc16f1f3fd290da90ad7f9a10f75;
mem[505] = 144'hf0f5fe4dfe37f4f90b0ffc3efe99fa43f2b0;
mem[506] = 144'h0a06fbde0f160b4ef214f0b5ff320b20018e;
mem[507] = 144'h0e91f4e8f801012e009af83f0c00f34706e1;
mem[508] = 144'hf02f02fc0ddb0998025b0a260ee208dcf239;
mem[509] = 144'hf043fde5f63df8670448f8e50894f4440c5d;
mem[510] = 144'hf04af4bd0ee3f3b7f934ffdbf6c2fdc8f4ef;
mem[511] = 144'h073af664fcc7f006f24b03d7fb4506ef0759;
mem[512] = 144'h0670fdfcf84df45bfb7e07f5f1c8f2c702c9;
mem[513] = 144'h09c90db7086d08df0d130c6af65008080e25;
mem[514] = 144'hf06cf4790d06ff95f71ef9dc0a60f73bf28b;
mem[515] = 144'hefe8056006fd0f8f046e0881fa040f1ff9a4;
mem[516] = 144'h02a0f9e108a3081df4650c5c0ea102affe88;
mem[517] = 144'hff3f05b4098b027df358f3c0fe21fdeaf03b;
mem[518] = 144'h070502560490f716084ff82af501f02cfc66;
mem[519] = 144'hf36f01d6ed17ee75f55c0392f60bef46f704;
mem[520] = 144'h061102c4006305f6f792f15a06d40ba0f65b;
mem[521] = 144'hfa960063f7af02c8ff8cf0d1f7c109ae0bff;
mem[522] = 144'h0baaf247f1e407090340fd30fad5033af115;
mem[523] = 144'hfde0069cfdd100b2ff12f51e010eff360a0b;
mem[524] = 144'h023f03f5f5a5fb26fd0ef49cf913fb2d0c10;
mem[525] = 144'hfbb0f1a5f949061a0280f939f7cdf261f34e;
mem[526] = 144'h04b1035df947f8c5095bf6caf9cf089e0125;
mem[527] = 144'h00c00ab50c4004a107b00386055ef26c0773;
mem[528] = 144'h009f02b4fb060634f32107bbfaa1fc01ff42;
mem[529] = 144'h058cf0c4f7c30cbaf09b02eafeccf6490456;
mem[530] = 144'h0cc4f3ad0676fb3bf9adf0d0f0580a6efd4a;
mem[531] = 144'hfd77f5fe040e0095f9cdfde309a90e34f882;
mem[532] = 144'h000bf468ee92ff43f3cc07d8fb0d0b35f17f;
mem[533] = 144'h059fefd1f1ee0b73f03df9be0c8fefc4f85f;
mem[534] = 144'h09430aa2033b098afeaa035008e5f5af01a1;
mem[535] = 144'hf5ed029508cdec69f52805c0fc55ff400b45;
mem[536] = 144'hfe510309fc6d0db4f9470a520605feb4062a;
mem[537] = 144'h0024082300fe0080f55cef1e0bd7fe370154;
mem[538] = 144'h0dcb0522f7cbf389f9830149fe36fe52f361;
mem[539] = 144'h0007f8a2fffef6e2fdedfdb40104f253f0d8;
mem[540] = 144'hff5a03b402fa0ef0f18f0e4ef591fadb0681;
mem[541] = 144'hf7e0049a047df94c00420a81f5d305e1ffee;
mem[542] = 144'hf9410d4af5a600900a650714fe37f3aaf62d;
mem[543] = 144'h0b6d0c580b6a0729f83409a20c7ef1ce00c5;
mem[544] = 144'h018c07570ce2007601250116042bf5e501a2;
mem[545] = 144'h013c0e8605c0f73e0631fc06f7f00acb0a4c;
mem[546] = 144'hfb7c0f650ca9f6d3f742f67107e3fa5e0f89;
mem[547] = 144'hf2cf07c201c3fc3800fbf2a80cd705b1ff59;
mem[548] = 144'hefb003c7ed5a0ee6f245f2b7f2edf433f6b9;
mem[549] = 144'h03aefd5bf5430d3a00c9f4360b75053601ee;
mem[550] = 144'h08a1096a0906fced0bbc06e7eecf0578f402;
mem[551] = 144'hfe62efca01a7fb49fbda00e3f70aed1bf9fa;
mem[552] = 144'h0305fa03023b0578fb16f00ef8d5017008db;
mem[553] = 144'hfc230d4ffc1e0287f3a0f42eeda60d3c0446;
mem[554] = 144'hfbc80e51f65bfeb3f73c070af209f57ffdc8;
mem[555] = 144'h07c50262f184fb5805e6f4ea05c00289fff8;
mem[556] = 144'h01d6fe3d05490afd03bdf6f30a0dfc4af4f3;
mem[557] = 144'h07f3012d03a3017cf24a0219f2890a02fed0;
mem[558] = 144'hf78504c5f08c0e46f514061d07670e3207ae;
mem[559] = 144'h0d13ff3ffc69fa4109d60d7d0dd3fc260897;
mem[560] = 144'hf830f97df0610152fd2ef8cb0c7b09e7f598;
mem[561] = 144'h0e2403aaf925f33cf647f9e5fc39047bfc40;
mem[562] = 144'hfd2f01530e55f752f0b2f225f34cffa00af6;
mem[563] = 144'h0b7706b6f512f17a09e2fded06ca090405da;
mem[564] = 144'h028ef93708e8f5160459004ef5cbee1409c1;
mem[565] = 144'hf8a4eee607c9fd0bf3b4f8ab026e05680179;
mem[566] = 144'hfac7f4560bf7fbc9024702e1ff41ff1dffd8;
mem[567] = 144'hf96604be099bf88507110190f857017a02eb;
mem[568] = 144'hfb91040f0dcf0d49f47cf2c20651f3d6020a;
mem[569] = 144'h0777fec3096efbd2ffad0530f3cd0de00c2f;
mem[570] = 144'h02f3ff59f886fc94fc8004b2091e0cfff566;
mem[571] = 144'hf59af750f5a204990779f1890b33f4710c14;
mem[572] = 144'h0b5700d3f0990ac705b0f2b9002f072b0492;
mem[573] = 144'hf2210724068407b3fb370b10fc1400b10a76;
mem[574] = 144'h0e25f81d082ff550f07affbe0bfaf2baf94c;
mem[575] = 144'hef18ffd1faecfc41fb380771fc3efb2c0c9d;
mem[576] = 144'h05fdf15cf43509cf0053f7a9058a070402c0;
mem[577] = 144'hfe8ef22f01f40a7f0a4b044c02cff2f9f542;
mem[578] = 144'h0267f2c40df90879f07bf000f18c0870f1ad;
mem[579] = 144'hfc19fa2305d10a72f4e20c18f046fb100cd0;
mem[580] = 144'hfb05ef80f2f3fd7af959fd210ae0050c048d;
mem[581] = 144'hf163054105150cf2f33c074c0b5efd6f04df;
mem[582] = 144'hf45cf15006cafe9df65603fdf87309cd0e0c;
mem[583] = 144'hef5d0862f7e3faecfa02ef81fd84f9e5f1ff;
mem[584] = 144'h09b00353f2dc08c8f139005ff6b00d76f489;
mem[585] = 144'hf88302eafb03f5060004088400aff2d208d7;
mem[586] = 144'hf67af3ef0a1f0334050df92ef65cefdefc32;
mem[587] = 144'h0bf50d91fe03f8a20961fbb00b7f0ccefe88;
mem[588] = 144'h03e10895026a0ee702eefe160b8f084d00aa;
mem[589] = 144'hf3baf98702350a4803c9044afb93fd2700b6;
mem[590] = 144'h0c300c07f8580f27fe93ff75f392f58b0ea7;
mem[591] = 144'h074d02970845f9dff33805150fb108920edc;
mem[592] = 144'hf4e60a96fc6009640c4ef90f05e60591f4eb;
mem[593] = 144'hff77f67d0409fd95f6f1075ef1670261078b;
mem[594] = 144'hf5f2f8310fe5fcac090f0457f5f1079b0747;
mem[595] = 144'hfc4ff6c2f5660480f8dafd770748f424f9df;
mem[596] = 144'hf04dfda40d9503d3f28d0e46f14ef466fbd0;
mem[597] = 144'h03e007effe490139fb770879f985f87108a6;
mem[598] = 144'hf46e0b7d014ef84709bcf8c9f95ff4e30c69;
mem[599] = 144'hfec2047300590124efc2fab5076c00b6f49d;
mem[600] = 144'hf99c011cf18cf7830dd7f463f934efdcf4d6;
mem[601] = 144'h0e31fbcd0589f574f3d004230a2502fb043b;
mem[602] = 144'h023a08bdfa580df3f140f7ebf4b5f590f64b;
mem[603] = 144'hfc80f451fb45084d0d49fe07f782fad80f2b;
mem[604] = 144'h0cad0a0d02bcf2420281f8580ed3fe25f3fe;
mem[605] = 144'h0c2e0cef0236f987f2abf92801310942f6cd;
mem[606] = 144'h06060562ff8bf6d60c75015e0969fc6c09f6;
mem[607] = 144'h0a01fcd40862fe84f0130e720b8e0b280383;
mem[608] = 144'hf008fbca0ae6000ff4c70ed106430d3ffe41;
mem[609] = 144'hf8c4fb82fcc20744f33007690c5e0ed30bed;
mem[610] = 144'hf0b5f6b6fcb30a53f09809b0ff21045af3ad;
mem[611] = 144'hf4e206a40c97fbc0f1770508fac50909f731;
mem[612] = 144'h0398f8c60371058df70908bff1b105720d3a;
mem[613] = 144'hfe0b0d1c0cb50ded0fd40fca08a9f48cfc22;
mem[614] = 144'hfb8ffd6f063b02d7f56e093b04d80b09fd59;
mem[615] = 144'hfd8b0bb5f7aff862f4d5f11afe7ff41a0207;
mem[616] = 144'hfec1f62d0bb5f0160095f814f9faf64afb27;
mem[617] = 144'h0d12fdb6ff03fabff13e07c5f52b0ab5faf8;
mem[618] = 144'hf5dcfb1ff717020700af051ffba60faafb3b;
mem[619] = 144'hf1f2ffe306e3f49bfec7fad6f736f9890720;
mem[620] = 144'hf964071bf5d0fdac06e5fd4cf119060ffdae;
mem[621] = 144'h05a2f71203b70daffd05fdd4f44105c2f0c7;
mem[622] = 144'hf060fd050ea60362f9d7f1b1f20a050ef726;
mem[623] = 144'hf3ca0a360121f416fab5f33f0009f6aa05cf;
mem[624] = 144'h01eb0513f6cef8d7fddff75a09920a3d012f;
mem[625] = 144'h047afd6ef7be0df903d00e6e0b4a0ad8fb3f;
mem[626] = 144'h050dfa11051e00cc0ce0fc9bf04df7f8ff88;
mem[627] = 144'h0ae3fc32f13d05e408dafe1509070409f313;
mem[628] = 144'hf3f1f9bcf7ac0d160a900d86f794f1610006;
mem[629] = 144'hf3d7fa77fc5aef31fa3b0b01fa3dff00f1ab;
mem[630] = 144'hfee9f42d01370eb40cf1f8abfdf2f90cfe2c;
mem[631] = 144'hf77aff87ff5aef7af91306f00ca7f0d80095;
mem[632] = 144'h0549008905e60106f8770c1ef5ebf548063f;
mem[633] = 144'h0d64f8a7f71104dafe530590f146084d078e;
mem[634] = 144'h05ebfbcbf51d0361f0ffef930178091d0b64;
mem[635] = 144'h022607c10a4f022f0ebafd0cf359fe070652;
mem[636] = 144'h0479f647feb1ffc7f97def94fb470cf10ce9;
mem[637] = 144'hfb0cf4d9f80e0268091b0209f61df65200ae;
mem[638] = 144'hff2f02ce011bf4b30fb90addfc4901daf67d;
mem[639] = 144'h031c04e5f1b7f55900f705ed024cfc75f9c4;
mem[640] = 144'h01700ca60de5f3d1f1df01270521017cfebf;
mem[641] = 144'hfcf1080f0dd2f97cf352f170f29607eef5b2;
mem[642] = 144'hfead0ceb0a55f349f648f8680b76077f0bcb;
mem[643] = 144'h0b820da8f9f3f8b00943f345f4e90f76fa4a;
mem[644] = 144'hf974f0eb05c30cfc090af739fdc4f05cf4cf;
mem[645] = 144'hf1ff010a048dfd720ca2f624f96ffb1ffd52;
mem[646] = 144'hff85f6f1fce20c0e08a00e6a03a30269fa25;
mem[647] = 144'h0ae40e9cf545ff3002fcf48efad60deffbf3;
mem[648] = 144'hf2d6026c0b0b0f94fd0406b2f8750eebefdf;
mem[649] = 144'h03f504f3057ef2510519fa84f682feb000a0;
mem[650] = 144'h0744f579f9d405b5f14ff48ff9acf67405fb;
mem[651] = 144'hf93f0e390aa60e07021ff4f4f4e405cafbcc;
mem[652] = 144'h032df215f7940250f9e4ff6bff6efcd1f593;
mem[653] = 144'h0908fc6303d300bf05ba0c6d0cf9fb700427;
mem[654] = 144'hfc5cfa0af37b0b1bf4e1fb1efa51fd620e0f;
mem[655] = 144'hf3640bf8f7d80d2e0830f9f1f08d00eafe53;
mem[656] = 144'h014cf89b0f050c5dfc07f664008ef07f0aaf;
mem[657] = 144'hf8b40d0afe54f9fd0970fcf8f54906480fbf;
mem[658] = 144'hf65d00a603eaf1820373f911ff26faddf088;
mem[659] = 144'hf1c703f60af4f410fb93f9f1035107adf0a8;
mem[660] = 144'hf662ff8aff9cf196f436ef9903b4099004fa;
mem[661] = 144'h073c03620e0a0284fe2ff5e7089907ea0854;
mem[662] = 144'hfcdcf96ff5300e550c8dfc5dfbaf0eb2f2c2;
mem[663] = 144'hfe75043f010e086ffa47f4f305390168ffb0;
mem[664] = 144'hf30bf58b01f20265f69ffb74f133028ff3e0;
mem[665] = 144'hf5ea0271f7ee001ff04a07abf3c0f4a1f52a;
mem[666] = 144'h01a1f405fb64f7eaffe50706feb00aea067f;
mem[667] = 144'h033cf7990866f24dfae6f4420c68f0ee089d;
mem[668] = 144'hfbc20436f1abf846f6900c8c09610749f5e8;
mem[669] = 144'hf5dbfdc00485f6250903f2b8076b0a57ff36;
mem[670] = 144'hfa8f017e062cfa56f683f9a4073cf293f19f;
mem[671] = 144'h043c0d2b049f0b3905f402c90ab6f2890925;
mem[672] = 144'h06250febfc010f0a0717fde1fa9cf3040fe0;
mem[673] = 144'h032203f700e801970cd9f007f037f7b50ea0;
mem[674] = 144'hf648f531066a0e0900b406d6f4ccf9b00a34;
mem[675] = 144'hf9a7f29bf37ef98bf9a2f8ebf3ea0ea9fa56;
mem[676] = 144'hffecfaf7033d0450fc47f642f76907410883;
mem[677] = 144'hf4ccf4f6f92908b3f7d70d31ffb9f39df913;
mem[678] = 144'hf272082af7240041f698fde7f88d0b29fda2;
mem[679] = 144'hf97f0c7ef20200790aceefbdeecbedf70980;
mem[680] = 144'h0a1c0f0c08a1f7d40031f0edfcf2fed80de2;
mem[681] = 144'h0ab8ff150a3308fb0ce0f68cfb46f23ff061;
mem[682] = 144'hf206fe7efa520124067d02e3009e0da5f0e9;
mem[683] = 144'h063905be0b4b018bf3ef0ceaf63d054ff302;
mem[684] = 144'hf45605c0024cf7f50cd3ef30017ef00d020c;
mem[685] = 144'hfb56000b0b08f7c7f0040881fd9f0cb60389;
mem[686] = 144'hf14d0e43fa3703160dcb0f47f34306e60a04;
mem[687] = 144'h008b0a1afefa037bfcfaf6a0f4a70b7d08e4;
mem[688] = 144'h0dae0ab20f830e29f30bf48d0de400780f1c;
mem[689] = 144'h09510e95045001aefa00068402e0f147f4fd;
mem[690] = 144'h0631f498ffaa03ab069df636f7daf4110915;
mem[691] = 144'h062d08fa07fff3940fbbf0250a3bf4a8f37a;
mem[692] = 144'h0b050fed03d5ff63f84b08fe0643f31a0b16;
mem[693] = 144'hf6da0f8207310f23f81f0553fb9e07df077b;
mem[694] = 144'h088afa08f3f50050fdfbfb5af4af0712fa11;
mem[695] = 144'hf2b6fe10fa430bb90c5709e008a1fa070476;
mem[696] = 144'hfc32fa0efb88036bfcfc0f300b20017e0fc2;
mem[697] = 144'h0729fe7e077cf1b5f8d7016f00f9f6c80603;
mem[698] = 144'hf1b80d04f8e5f48bff74f775f1b1f36f02be;
mem[699] = 144'h0db1f0840a6d0ba300b2f6ec0572076ef4a0;
mem[700] = 144'h012300a00a8208770b050b1e05c00b3af8e4;
mem[701] = 144'h09a10e4cf03701c4f6d6f17308dd058b04e7;
mem[702] = 144'h0dccfdedfc08fd9f008bfb9e0f600c98f060;
mem[703] = 144'h0ad30ce60c37ff9dfe49fe88082ef5bf02d4;
mem[704] = 144'h0e360952f3e8046b0559fc03f7e30e7a07de;
mem[705] = 144'h0f1108290560047ef90208f706a4fec90db9;
mem[706] = 144'h07eaf20c00480fbdfb4d0290f1d1f053f632;
mem[707] = 144'hf5180611ff1b0f6a0169f500f56b06ec02b7;
mem[708] = 144'hfd43008a0705f93303190e8b0129f683fea1;
mem[709] = 144'h022fefd107cf0adbf4d9f29c03ff0374f2f5;
mem[710] = 144'h002cf09ef66101be04c5f8b7007b057a0f9b;
mem[711] = 144'hfc7b04ff0715f89e0391f458f9b0fa3cfa7f;
mem[712] = 144'h0a8cf6470c550d79018105e7fb3a060cfb29;
mem[713] = 144'hf10dfe3301faf16705effccbf1a007cf0cb2;
mem[714] = 144'hff1cfc49f97403f30783fdcaf39bf4d801be;
mem[715] = 144'hf1c90d400b74f828f27a0cd20a83f3a4f302;
mem[716] = 144'h0d2f0ad8f91f0a11ff6308170c43f37c089d;
mem[717] = 144'hefda0ea70526ffd8ffa8fad20b840f990195;
mem[718] = 144'hffcb027af715fe83f3f003140ab908b0f2be;
mem[719] = 144'hf676fa5706e904b6022600100f99f2a0099a;
mem[720] = 144'h0ce705020859f2e6f97a0962005b0afaf666;
mem[721] = 144'h08bb00cbfe0b0317f03702120848f3b8fd96;
mem[722] = 144'h01620b5908f3ff410848f7ebf6910d990d36;
mem[723] = 144'hfac1f328f98c09ecf04a0bbaf574f8ee0c50;
mem[724] = 144'h02120bf0f14f07120541f705f125f25af2c7;
mem[725] = 144'h040ef61ff5c60fb301b1ff6df5f70cc0f54b;
mem[726] = 144'h0d6f0a7ef1f90b290fc40e430075096dfde0;
mem[727] = 144'hfe8b0316f9a7f5ae099d081ef745f544f844;
mem[728] = 144'hf06ef861f40601bef89ffe360d9af417fa77;
mem[729] = 144'hfcfbff51057ef34ef42600a30928fab3f418;
mem[730] = 144'hf9010e51fc39010b0deefe2cf5f401520ebc;
mem[731] = 144'h05310cdef6acf8f902600cf5f937fd580350;
mem[732] = 144'h080b0d5ff72a0ac2f8100375fba8f409f737;
mem[733] = 144'hf8adfed60eebf2ea00500793fbf1feef0390;
mem[734] = 144'hf88a04adfca20c6bfbbafde0093202cd06ec;
mem[735] = 144'hfc7df5730e5efb90f0bf06ec0637f3ee0c0d;
mem[736] = 144'h0343015e028af264032509f907a90de8f126;
mem[737] = 144'h02ff0b0ff562f528ffddf0bef6c1f505f715;
mem[738] = 144'h00d20f2ef14b0f71002d0df2fee50d1e05e0;
mem[739] = 144'hfb27f61b02ebfef70b590738f46f02ea0c8b;
mem[740] = 144'hf3c0096609500027f2570bfbf4de0b10f40c;
mem[741] = 144'hf6acfe9a01ba0453f5d0f47f06f0067c0d2a;
mem[742] = 144'h01550f780c390ac6f18bf9ca013b0971fcad;
mem[743] = 144'hf639fbbbf108062f0a770dff03d0fec8f85c;
mem[744] = 144'h0ed009fd0240fab4090f09a80539fb5b0386;
mem[745] = 144'h03490e410ad4f0740d1c0e24ff72f4cc067b;
mem[746] = 144'h0b020e680b69f21e0e51089b03740af90d3c;
mem[747] = 144'hfe6efa3d0b6605b10f23fefb0c010597f7e0;
mem[748] = 144'h08a5f20ff13df33306d4efc90625f9faf3ed;
mem[749] = 144'h0c94ffcffe5ffce709ca0b6bf59e04b10260;
mem[750] = 144'h0618fc920cc1f068f8a30615fefff74f0f71;
mem[751] = 144'h05a0f6af0f450943f00300ecf1c503e509b1;
mem[752] = 144'h0da3fc5f03e0f5d6f4db0cebf8220f26f609;
mem[753] = 144'hfe5e0a1c0638fd5f0fa1f03d0eeafd6ef45d;
mem[754] = 144'hfd030dba0cd5024e08810210fec0fc3a0c6d;
mem[755] = 144'hfaee0ddff6cbfc2c0300f23cfde8fefa0122;
mem[756] = 144'h029afa62fc9d05acfc900e4c02c3f0c90247;
mem[757] = 144'hfe4901d2f1f4f501f3260c04f869f3c20939;
mem[758] = 144'hf72c0f560761f41cf930f842fefdfb32fca1;
mem[759] = 144'hf227f4380750fb2cfb42fbfb0edbf4c90c56;
mem[760] = 144'hf3620c100712fdf4f1040d21020bf91b0049;
mem[761] = 144'hfe470fd8f19ef9260730ff96fbbdfe70feb8;
mem[762] = 144'h05090f950688f0eb03ad0f8c0f8bfee70846;
mem[763] = 144'h0ecf0beaf0fcf5420e4ffd1703ddfe6207c9;
mem[764] = 144'h08bcfbfef35206fb0a43f0fb08450c3d08a8;
mem[765] = 144'h0cac0ac9f7ee05590b9f0fd503b30a070a87;
mem[766] = 144'hfd460bc90d8efdbd09f70144f07b04430293;
mem[767] = 144'h0da8064df6090ccdff0bf4ee036103070fc2;
mem[768] = 144'hf3be0a4bffadf103fdf6014a0b0ffbeb027b;
mem[769] = 144'hf4cff4240d95fbcf07920fa0ff7a054ef853;
mem[770] = 144'h01d2fd1a076cf770fb990c25fb3b067106cf;
mem[771] = 144'h0c4ff5ad05c805d60b01f4510bda02000816;
mem[772] = 144'h042ef734f4330994f6aaf529ffa4f764034c;
mem[773] = 144'h05e7f75a0533f049f8cb0b53f6c90b160823;
mem[774] = 144'h056802d8f3bdf7e8f4def1580457f091f527;
mem[775] = 144'h05bb03730163f9ddfb0107ff00e5092cf2c3;
mem[776] = 144'h0660042106c807120599f652f50b0bfe01bc;
mem[777] = 144'h0412f81bf0c3f65b075af2b00306f7caf76f;
mem[778] = 144'h0ee2ffda07cef6130dec07020b75001df79c;
mem[779] = 144'hf284028df172fa97f3150f45ff40fb51fac3;
mem[780] = 144'hf9f5f4f0075f08bc0ee5f762f719ffb3ef6b;
mem[781] = 144'hf2a7f5a9f44df72af26ef83109e902940093;
mem[782] = 144'h0d05072e026e0dca024b02edf69bf294f1a1;
mem[783] = 144'hfbc3023af5b505baf345f3d60f7b0c4e023c;
mem[784] = 144'hfae60304f70b0732f0670a290137fa44041a;
mem[785] = 144'hf69e083afbc2f290f9e9f670f1fb0f1a015e;
mem[786] = 144'h07600cd903b4f3be0d990fc4fe1c0583ff84;
mem[787] = 144'hf4d4f0d5f910f33a08a60dc2ffad0cfafd08;
mem[788] = 144'h09f9f80f0c2f05cd0dfe034a0f93031f05e4;
mem[789] = 144'hefe70f2d04f30dcbf6d104520009f1680b6b;
mem[790] = 144'hf8950242f60cfaaa0d4ef94afbff018afd2e;
mem[791] = 144'hf535ffc0ef1bf706f03df3520984feb60ab1;
mem[792] = 144'h0e820cf0066bf70d0bb3027cff6ef4f30cb3;
mem[793] = 144'hf7d308230bbd0c5ffc7ffd3ffd04ff3507c9;
mem[794] = 144'h06f8f0e3f79cf6b8ff920ad6f9ac0fd3067f;
mem[795] = 144'h09780507012af77dfd7306e603ed02a30846;
mem[796] = 144'hf18ff3220691fdd202900acdffd502450be7;
mem[797] = 144'hf27bf81d01b4f65906cc076cfd5bf1850519;
mem[798] = 144'hf7eff047f206fc83fd7d0958f97df80904d1;
mem[799] = 144'h0bebf18afb5e034c0eb800f1f9d0fedaffce;
mem[800] = 144'hf0e608cef49cf49cf74b069b0d18090efbac;
mem[801] = 144'h059303130464f78f02c5098af538f8c1f29d;
mem[802] = 144'hf95eff7e082af42a0ccf0e46fa8af4150aa9;
mem[803] = 144'hf461004ef5c6f089f2a30b800173fc8df042;
mem[804] = 144'hfe64054b0ab7f363f93f07fa0d91fdc0fb09;
mem[805] = 144'hff65fce8f3c2f2b302a9efa408a1ef4d0bda;
mem[806] = 144'h0a7bfae8fc8a072bf319f315f600f7480023;
mem[807] = 144'hf605f2c103b0f524fcd0062efa16fd24fb4c;
mem[808] = 144'h0328fe790796f4330c1e0cc60c93fbcc041d;
mem[809] = 144'hf4070a5aefb6f94df65c0ab602d40a15ff53;
mem[810] = 144'hfa0e0b42f403fdda019ff3c5f5d2f5f0f535;
mem[811] = 144'hf68c05baffa408cc0516f726ff8dfe490a98;
mem[812] = 144'h0c7f02d8fd2cf2d507e9fd2af78d0e85f21f;
mem[813] = 144'hf188021bf9a604f30b4ef546ff38f14506df;
mem[814] = 144'hfa56fec6f74f069008f706f205630455fa99;
mem[815] = 144'hf450f679027707330c9ffeaff7280491f0d4;
mem[816] = 144'h010c0f94044d0459f86df15cfb34f6ca045c;
mem[817] = 144'h0e36fc790c460fd108fafb5cfab500ee0309;
mem[818] = 144'h091bff07f91a07bd01a7ff4e024df66ef2e7;
mem[819] = 144'h0d40eef4f953f606fbb4f940f1c0f210f600;
mem[820] = 144'hf49b0d8d09280e77f8b2f8c0071e05e5f367;
mem[821] = 144'h0032f0dd0b3d0107fe470d8bfc2ff8410c59;
mem[822] = 144'hf8610b6f06e0057df1870739f0befb30f8be;
mem[823] = 144'h004feef1061606dc03bdfd3bfa8ef6aff727;
mem[824] = 144'hfa8701e9ff32f40408c4f85905520601084f;
mem[825] = 144'hefb1f5d6fa2c01a6f75e0d2cf0bffcab0384;
mem[826] = 144'h0efaeff6f9850016f96ef5fc0d10f894fb5f;
mem[827] = 144'hf7c0059dfb4ffda50983f61808a8064707dc;
mem[828] = 144'hf0720623f2aa084bf3e00791ef9a0000ef3f;
mem[829] = 144'h0e24fe380b5f09bb0ac700f106a20ebaf2cc;
mem[830] = 144'hf9a1037c02fefb560997f269089ff87df63f;
mem[831] = 144'h01530b6c0d730808004af929f5a30083094a;
mem[832] = 144'h076a091709a909460059f4a60dea0eab0c83;
mem[833] = 144'h03fb0ab3ff640d17f382fea30c0c0db2f0df;
mem[834] = 144'hf26cf55ef699f46c00a9f3fe0fc10ce3f0d0;
mem[835] = 144'hfdfc01c80d7ef8230eadfe2efd960817f6f3;
mem[836] = 144'h0c1003720262fa91f29df4b1f6b9f555f96e;
mem[837] = 144'hefb305c6f50008000d2f040a037bfc0afc5c;
mem[838] = 144'h043a0a2cfbd1fa37042af8040c66fd3604ab;
mem[839] = 144'h064c05210a680a940a13f1b9ff02f8ecee87;
mem[840] = 144'h08520728fb4706b0043afada0b87fc3cf827;
mem[841] = 144'hf0010f4bf22bfe0e0910f178f5a6099805d1;
mem[842] = 144'h015808140aa5f08f0ad507a9f844fbe0f2ab;
mem[843] = 144'hf3b1ff68fa02fc0a0b4705df0ea1efe2fa47;
mem[844] = 144'hf79100bdfc520e340597fb3a0b63fe7f08dd;
mem[845] = 144'hff9109fd06aef2de0079f352f42e0965f0ac;
mem[846] = 144'h0c14f3d5070f0f930779021efd2c0eb8f36e;
mem[847] = 144'h0deefb49efeb0895f6cb0a73fe6808740c26;
mem[848] = 144'hf5980b430566021cf6ddf7570d9f0dabf810;
mem[849] = 144'h0c11f11703f1094e0286f339f11ef51ffe76;
mem[850] = 144'hff14f2a604def5fbf5b8f20c06f70c89fabe;
mem[851] = 144'h0646fdc704fc0f13ff6c05d805c7fb8301ad;
mem[852] = 144'hfb7e0a3efcf3f9ed03dc058a068100e2068f;
mem[853] = 144'hfd85f6c40076005afccdf1adf4adf832f855;
mem[854] = 144'h0009f88ef8d8fb21fdff09f6f10e03fb03be;
mem[855] = 144'h0881f28200530357fe1303eff780fd110928;
mem[856] = 144'hfe60f302087d04e300750d7f0e9f09fff52a;
mem[857] = 144'hf98707f604a1052ef4ff08040b71ef6cf947;
mem[858] = 144'h00bef846fecd061e002cfc600517f117f6af;
mem[859] = 144'hfc5cf81dfc68045807c3f22e09be00df09b3;
mem[860] = 144'hf886067bfeca07cd098c05600436fcebfde3;
mem[861] = 144'h0cd7f145f01fef730b420f57ff86035cff97;
mem[862] = 144'hfc90f0830d43f3bafa25fff9f6b206cf011a;
mem[863] = 144'hf0a205820cf10b44072cf327f62ef22d0142;
mem[864] = 144'hfd69ff6aff14fc0afaf3f7b402bdfba8f91e;
mem[865] = 144'hf577f22ffe9cf4530b9b086afafc08b5fa6b;
mem[866] = 144'hfcbe04420db3fcaf037afc5ffb8bfc15ff94;
mem[867] = 144'hf111094906cff5c7fb6cfc670e0bfe04f12a;
mem[868] = 144'h09e40846ff3104e6fe7000bf03fdfca8f407;
mem[869] = 144'hf8e7f8a2f04ffe10023af78a03fb03a106ea;
mem[870] = 144'h05cafe30f311fa0bfbc40715f8480a340621;
mem[871] = 144'hfbaa05f6ef230406f5c3fc70ff12ec660877;
mem[872] = 144'hf770f950f179f032f7e50005fcb00a9f09c7;
mem[873] = 144'hfcadfddf0ac50be6f97101f4ff56ef58f1c3;
mem[874] = 144'h09f80c20f662f48ffc7cfd41f8baf34ef74f;
mem[875] = 144'h0906f5b6f74e06830a450bc2fd5400c5fd96;
mem[876] = 144'hf0a90e1ffeb4f23b0742f68b0b79f5d2fedd;
mem[877] = 144'hfa06fb3c03a0f247f82c0891f5a7f790fc3b;
mem[878] = 144'hf465f271febdfa00fca9ffdcf1c8fb33f026;
mem[879] = 144'hfb76ffe4f521fcbe0b51f3fcf873f738f603;
mem[880] = 144'hf2e00bea0e330a4907e8f568f338fb01f3fb;
mem[881] = 144'h059e0e00f342019c0605fe5c0444f3150e19;
mem[882] = 144'h0d26f9f309bffabd074801d10253f801f736;
mem[883] = 144'hf5c601fd0e45f168010f0033fa9ff8b7fd24;
mem[884] = 144'hffec0081000bf481f81afdf502e00da706f5;
mem[885] = 144'hf9fdf76708e105def1a807b0f880f70f0d22;
mem[886] = 144'hff19f1a6091bfeb50942f783f1920b7af7da;
mem[887] = 144'hfd8af06af81ef630f54700f7faedf6fd0b21;
mem[888] = 144'hf58dff71fd41057ef2a503e50902060ff0e4;
mem[889] = 144'h0b1c04dcf7e2f4550ceb0c6af6ee03aef0e3;
mem[890] = 144'hfd68fe4e01940f7404e9ff69f3feff73f79e;
mem[891] = 144'hf02eff24047c0d3107d2fba5f8c90785003d;
mem[892] = 144'h0985f7e6f953f156f030f82e0d2304d7f00a;
mem[893] = 144'hf046f2bffc5ff7e50744ff09f5b7efcbff37;
mem[894] = 144'hf5530277f54908affbec0babfa73f8e7f22a;
mem[895] = 144'h008af969f0a2fc02f6800020fcc1fe9c00d3;
mem[896] = 144'hf9affaaa02edf9c1fd3cf785fbbd062800e5;
mem[897] = 144'hf9e1fc93f394f1b9f7c6f9810a7c0c41f9ad;
mem[898] = 144'hfdb2feecfb36fead0c070d84fc2b034901c0;
mem[899] = 144'h00fff081fd3af2b80ef40df0f32803050260;
mem[900] = 144'hef41f67205ebf8e1071cfdba0a31f946fbf0;
mem[901] = 144'hfcfaf1b201f9f7f5efe0f5200e7d0e5ff7dc;
mem[902] = 144'hf6a8f007003c0bd8f1db05e2f2cc0e29ff97;
mem[903] = 144'hfde3f65afff60cc708eb0615f1bf03a4f72a;
mem[904] = 144'hf53ff3820f44ef5401ba095c0267f93af300;
mem[905] = 144'h0380f32800a600b10d740a31001909620726;
mem[906] = 144'h0fcbfb2d08130eadf1ac0b65f293f9b5038f;
mem[907] = 144'h09680f96f4dff9dd021504c909520c60f48c;
mem[908] = 144'hfcfa0552f456f70ff64a0748fcd20c8f081b;
mem[909] = 144'h0a290de2f854fbb20ce60232fd58f32afed9;
mem[910] = 144'hf2b009f3fb070d34fd46f0b40bb0f054f8dc;
mem[911] = 144'hf4bafe02fe6b0b7efd04f484fbcdfee000c9;
mem[912] = 144'h08f3f690f741fa38f1c7f8cdf8d206ee0a43;
mem[913] = 144'hf05900cdf36d05a6faf3fb5bf16300b2fdb4;
mem[914] = 144'h0e3ef6c1f8a5f349ff250de4fbe8040305cb;
mem[915] = 144'hf98a0575f978fb4bfe18ffb1f82f0b050ad9;
mem[916] = 144'h00e4fb34fb31050f0e13f35b012af5e8f050;
mem[917] = 144'hfbc201abfc7ffeb8f3ecf060fe01050dfb77;
mem[918] = 144'hfcd40abd03460e59f207f2f50e970c7dfa45;
mem[919] = 144'h0681f161f46d0ab3feaff5beffc5f206f88d;
mem[920] = 144'hf4520777024d09440ccd0c0e04880aecf906;
mem[921] = 144'h06e1f46ffb7f0623fa68f3f00d75f965ff02;
mem[922] = 144'hf4f6062f06fafd31fff8067efde3f70af30f;
mem[923] = 144'hfc74fe70faeafbee031efe8af146f8060d9a;
mem[924] = 144'hf055022e0e1cefb7fc20f2e9009bf85bfdfe;
mem[925] = 144'h0ac00802f72b0cadf7a10e90fc9cf34dfd78;
mem[926] = 144'hf2800be609f7f022f0ae0f89039809340f7f;
mem[927] = 144'hf4ba031a0dadf128ffdff75d0c5cf9b3f4e1;
mem[928] = 144'h011cffbd05dd091efc750e66f8780992f991;
mem[929] = 144'h09f30ca7fe350a50016eff52090d0f08051a;
mem[930] = 144'hfcf0f00b07d3f572080b0a5efd93f0a10ab7;
mem[931] = 144'h0d67f3840b340a750b0a095d0efa04090573;
mem[932] = 144'h095100acf78101300e6fef100b8f01ab04ac;
mem[933] = 144'h0310f79403c10ac9f3daf33afa1e0469f7dc;
mem[934] = 144'hf852f2cdf16901d20df406550080f3780496;
mem[935] = 144'hf7cf0baf05f4f5f60cd90d4ff20b0d32f7ae;
mem[936] = 144'h00e500df07b301cffb47fc7af1ac0b520175;
mem[937] = 144'h06b40862fcd2f890eef506abf6bf07ad0768;
mem[938] = 144'h02cd0b6d0740f7d409f4f161f9f2f0e1f2b7;
mem[939] = 144'h0e620d7c0b3c0ca4f3a9fb71f549086ffeae;
mem[940] = 144'hf6bc0e58000b0257089bfba6f908efa805eb;
mem[941] = 144'h04790089ff04f072f67807640797032b0b9e;
mem[942] = 144'hf5190adef48bff07077df727073e0f57fc6b;
mem[943] = 144'h0db6fe8bf5030c24042f0c480eabefc6faa9;
mem[944] = 144'h0893f0f9fa42001eff2dfb13f73d02fd0932;
mem[945] = 144'hfdb8fad50def0d2af228fdc8f19d081cfc28;
mem[946] = 144'hf7bd098607220486f5cbf5df07c70a3b0caa;
mem[947] = 144'h02b30deafc7cf0c0f463075c0a97ffbc09d1;
mem[948] = 144'hf6b9f1050513f8f30a4c0ca3f04aff150410;
mem[949] = 144'h067af0ddfb8602a3ff0cfaf8028108fbfee8;
mem[950] = 144'hfab40001fd4b0e18024b046e0b3306c70f4c;
mem[951] = 144'h0917ef3904ad05360c90fd590ce70e85fb76;
mem[952] = 144'hefabf3fdfbd70c04f8d1fe57fb45f7f0fe10;
mem[953] = 144'h086601220bd906bef39bf5acf020f7d10cbc;
mem[954] = 144'h0202052807ecff5e0b62ff22f7aaf062f641;
mem[955] = 144'h0e22fe8e0d2706b4fa88012afc3af3fcf867;
mem[956] = 144'h0122fa2e0771048ff604f8a20608038bf2c5;
mem[957] = 144'h029807b1faf70fd30282fa000267f58c0786;
mem[958] = 144'h0d3c023c080409a3026d0cc6f879f26702e4;
mem[959] = 144'h04adfeabfaeb0f660d6ffb05f950099ff13b;
mem[960] = 144'h04680a6f07f5f8580a50f965f004f31bfdfa;
mem[961] = 144'hf2b904fa0430f4b5fd21065cf97006eff437;
mem[962] = 144'h0beafbc70b6a0934f0aefc94fb850093fe00;
mem[963] = 144'hf38ef08006e5f3baf288f46107970ca7f1e7;
mem[964] = 144'h0434f9e9f02e0efff55af4b70249f8750636;
mem[965] = 144'hf71604080f900f17fc9b05920bcbf19d0e2d;
mem[966] = 144'h05c70a5f0a950a520f180bd3036b0417089e;
mem[967] = 144'h058ef342ffb3f5fafbe7fc7ff929f3a3f3d6;
mem[968] = 144'hf147f173017cf497f6bbfeebfe690dde0d6d;
mem[969] = 144'hf9270b320b58034502cdffebfd4ffad60923;
mem[970] = 144'hf8f603e2fe470e1309370ae70d4efa3207ad;
mem[971] = 144'h0efcfa040f8e0e130ece03270a21f0ff0955;
mem[972] = 144'h0ce40de9ffc8013afffa04e30e15f0750e58;
mem[973] = 144'h07fcfe66f8ecfb4e0031f2f60d8f012f0c44;
mem[974] = 144'hf73c0dba08bb073f0c6bfef3f414fef302c3;
mem[975] = 144'hf35a024efea9f1f4faa1011cf43af91e0436;
mem[976] = 144'h0c7ff8650fea076ff9b6fcec0c8e01dd019c;
mem[977] = 144'h0d8107310d9ef9c1f7960558f894f00bf300;
mem[978] = 144'hffcdf07c0d66fbeaf4200d34040b0d1afcc9;
mem[979] = 144'hf7c1061103f2f53bfa4508b60824faef01e6;
mem[980] = 144'h060008ddfb7b01fb07f509bef877fc6c08fa;
mem[981] = 144'h0584027605fb0d6e07edf1f7093af70ff290;
mem[982] = 144'h0675043afc67f82ef58afb4a0840f1eafc53;
mem[983] = 144'heeff0ee00363055cf154fef20615fc74f41b;
mem[984] = 144'h0b1af3220ca500e2f157fc67fa3bf0210f84;
mem[985] = 144'h0f38f3ed0cca0be4f8b5fdedf0000d6ff2c1;
mem[986] = 144'h0c36fecdf6faf61108360dc1f5a2ffaa0750;
mem[987] = 144'hf5e30a18fa8bfb1bffddf4be076ffcaff1cf;
mem[988] = 144'hf03af0e20b59f71afb2bff22053f0bdcf725;
mem[989] = 144'h086fefcdfcb007d0ffe7f627f96601ed018e;
mem[990] = 144'h0845ff5afe050844fa7502190ee8f128faab;
mem[991] = 144'h047cfd330a51fa1bf29802bf0f4d04ec0edf;
mem[992] = 144'hf1c30591f89ef5340a3af983fe78f1560f85;
mem[993] = 144'hfc65f6d6f1d108f4ff89effc0d22f65bf999;
mem[994] = 144'hfd6206e1f89bf9cc0b6d01130b4af3cbfe15;
mem[995] = 144'hf3c206dc0a5a0dc9f15ceee90dceef05f288;
mem[996] = 144'hf9bbfc11072406dbfd76fe0405b6fd1b0480;
mem[997] = 144'hf528f46ef5500d9201acfef504a2fe67004c;
mem[998] = 144'h024a0335fccdfa660d94f47af23b0811fe29;
mem[999] = 144'hf2d3f7520af0f8a50b5fef7007cc02cd07fe;
mem[1000] = 144'h005bf1690c4bfb6d0b9709e0f09bf3bd0264;
mem[1001] = 144'h0e6cf191f9a5fb8308960df70070fe130d00;
mem[1002] = 144'h005ef29b0d8bf211f6940c5dffe70877fe3d;
mem[1003] = 144'h06810289f1c502f2fa0709a803b2f53ef4df;
mem[1004] = 144'h0a78f0eb022bf58dfc0ef42d0927f86f00e4;
mem[1005] = 144'h0cf7004a0d43fc45faabff2004edf6be01fb;
mem[1006] = 144'hffc90bbff2f6fca3044c0ac8fc690017047d;
mem[1007] = 144'hfda0f771f504014ffb37f90a08b6f437ffc9;
mem[1008] = 144'hf59d09660dd10d790218083a0282083e0612;
mem[1009] = 144'h029401acf9ceff9709cbf283035af8500a5c;
mem[1010] = 144'h01acf6fe06050cb9097efe72f3d70e46f9e8;
mem[1011] = 144'h05770579fbe50fde014b06c00babf125069d;
mem[1012] = 144'hf013f66cfa2d0c22f3eaf9aff5cc07fef860;
mem[1013] = 144'hfd0004db0980014df629f34c0e890a53f8d5;
mem[1014] = 144'hf1960562f8f0f5570494f58bfcb3f9dc019b;
mem[1015] = 144'h02d2ed62ec130397f706f970ee89fede03c6;
mem[1016] = 144'hfc32fb65fd78fb10f4eef9d7fc2ef4c808be;
mem[1017] = 144'h0cecf50c08b7f637f37d009901c8f320edac;
mem[1018] = 144'hfb1c05db0fc2f67e0ab60e2c030ffa960b30;
mem[1019] = 144'hf837f387f18dff4401acf8a6f47309fd045f;
mem[1020] = 144'h0c88f2b001b208b4f927f6450ba0f08df31e;
mem[1021] = 144'hfb79fc4af4ec0c0b0318f04bfea8f794fb2f;
mem[1022] = 144'h0cbf067ffc6c09750151006bf7730656f4f9;
mem[1023] = 144'h08450c360e11f630f63ef57bf517f1b6086d;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule