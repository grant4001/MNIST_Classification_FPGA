`timescale 1ns/1ns

module wt_fc1_mem1 #(parameter ADDR_WIDTH = 10, DATA_WIDTH = 144, DEPTH = 1024) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'hf479f435fabe0745f8edfee00320f09204d3;
mem[1] = 144'h07a80549f498fa76046ef9bd0f1c0038f4c4;
mem[2] = 144'hfc3bf147f490f279f518023a0c0cfe130c6a;
mem[3] = 144'hf59c0c3bf1b10a63086b0811f8810c100938;
mem[4] = 144'h0a15fe6e0d33f1a3001b036908a302750c82;
mem[5] = 144'hf56e053106260c9a02fcfeb4f0aaf7b40715;
mem[6] = 144'h03bdf22c024efceef2f80ec9082e029209f5;
mem[7] = 144'hff9bfe240eb2f90ef56406100723f3ac07d3;
mem[8] = 144'hf77f0f5c012d0f65f7f8f019fe9b0226f414;
mem[9] = 144'h090b07daf1260a22fd0bf1c3f0b7fdfe04cf;
mem[10] = 144'hfd960f31f84003ee0aea0cb10b91f49df9c0;
mem[11] = 144'hfda9faae0728f2b5f5c8f3c6f68d0f670de1;
mem[12] = 144'h0ed804e1f0f8f1a10b38083c01ab0e2103da;
mem[13] = 144'h0261f5eef1900e6afb540cf0f8c00ed6f35e;
mem[14] = 144'h00bd0fbefffcf5bf0202fdbb0b82f17c0f58;
mem[15] = 144'hfe6d0bd00f7ff135f00cfbfcf49af99afab6;
mem[16] = 144'hf287f20b0e8104d4f84df98af12af530f4ac;
mem[17] = 144'hf355ff730dcb03adf80e04cafda90b5100ce;
mem[18] = 144'hfe530b9800eb00d3f68303780e680883081a;
mem[19] = 144'h00d1031b0b120c2509db054b0e2ef1d4f3da;
mem[20] = 144'h0d970b69f61bf0e8f157f049fcd202d4ff27;
mem[21] = 144'hfdce0a0efa4e0d00fb4b048b0e2bf6860f1d;
mem[22] = 144'hf37308760e49063cfb840c40f05e06caf2fa;
mem[23] = 144'h0284fb4705210aeafa76fe0001520ee50a57;
mem[24] = 144'h04b4fa9d07b809dd083bf82b090cf09efdd4;
mem[25] = 144'hfee3f558f86afd8dfb8f0fd1fecb039ef6c4;
mem[26] = 144'h04de0612fb4cfe20fd72f9adf457f51007c2;
mem[27] = 144'h0da6f0ebf7ac05e0fc2700e6f2a505a5f408;
mem[28] = 144'h0afff9c303b2f50ff00904720be4081efba7;
mem[29] = 144'hf7c1004ef4ce0c5602f507cef95dfebf0d1b;
mem[30] = 144'h061503810691fc38f08e0f4802a4fa8aff47;
mem[31] = 144'hf813f50ef4dff95ff4e7fb1303860baa07e3;
mem[32] = 144'h0870f16808010507fee1f0b5efb6fdc30630;
mem[33] = 144'hff81fa1afd6f02d4fcd2f8200b15fe2ef8ea;
mem[34] = 144'hfa97faddf01df0e9f39ef966ff5c0ffe09aa;
mem[35] = 144'hfb8efe4e0e57f0bcf982fed1f05df46709ce;
mem[36] = 144'hf8e2fc53fa290bbc00c2ee6cf999ff98ec19;
mem[37] = 144'hee440b9dede7f450f191fec3fb7805fe0717;
mem[38] = 144'hefe1ff37f101f60aff62064cf994f33f00b3;
mem[39] = 144'heec0f713f09f0823f1bfe8d1feb4f120ff3e;
mem[40] = 144'hd9cfe6b505d8fcd0eadbfb24eeb5f3bd0ae1;
mem[41] = 144'h0bc107e60a0501d600e501a90745ee1e016e;
mem[42] = 144'hf286f7fbfbf7f513ee29f9c70721032a0af9;
mem[43] = 144'hf892067df65cf530ffd70a70fd6205540ef8;
mem[44] = 144'hf864f8d202110c25f3d7042a041c0d15024f;
mem[45] = 144'h0a5d059efc4efd5d0e7df9860571f4690202;
mem[46] = 144'h05f3ff02f3ad0f880681f9de0c680654fe30;
mem[47] = 144'h08ed02d004d3f2650019f764fe6904140663;
mem[48] = 144'hfbe4036afa9b0db1ffc9f859f98b081903f0;
mem[49] = 144'h09acf79bf1ac05e6f3c1f54b0ae8f81a06ac;
mem[50] = 144'hf496f37cfd99091e0e30fa47fdcaf82ffe18;
mem[51] = 144'h08f208b8f8c8f71eeef90b10ffa1f15506c8;
mem[52] = 144'he86bf74704fcf7d7ff23ecedff37ef3ef81e;
mem[53] = 144'hf6fc019303c1f891f435f1930780fd07fc0e;
mem[54] = 144'hff07f50e06fff172f3fc06c4f652096af533;
mem[55] = 144'h0784f460ef8a00c5fb68f066f28dfa3df269;
mem[56] = 144'he733feb0f2fffd8400faf12bfc92f1eafa3a;
mem[57] = 144'hfbb4f4d4f8dd0766fc370937080ff2c006f7;
mem[58] = 144'h0c98f577ff70f6cdedba03550235019e0f29;
mem[59] = 144'hff0f0725fec00297fd4f0a46f17af066ffaa;
mem[60] = 144'h0b4bf9900dcafbb3f874f02e025df83efb3a;
mem[61] = 144'hf28d01bff2d60645f7330bf9f059f8080a19;
mem[62] = 144'h04ccf5bd0126fe410a37f7a4fb850a23f7c9;
mem[63] = 144'hf8da08200c47ef01f1cef6def5de0894feb0;
mem[64] = 144'hfd06fc23042600fa0866f0d2f0ce04c2f15f;
mem[65] = 144'h09b50eb9058bf54a0ba5fa60078503600754;
mem[66] = 144'h09cb02f2f72df9db060502da03970c57f266;
mem[67] = 144'h054f095ff74909cf0b200331eed201520230;
mem[68] = 144'he231ef2eec73eeeaec78f37ce705fb06f451;
mem[69] = 144'h011ff8d7f2f3eea6ee02f249ef03edfa062a;
mem[70] = 144'hfc78f8b403aff65cf1f30956027dfecc03f0;
mem[71] = 144'hf49308570871f708fbddfaca019f07250b93;
mem[72] = 144'he55de737e75bf3b1ed16ee5afaf9f03deeef;
mem[73] = 144'h0bdaf657f75606aa0bb9fa27fe500a78f029;
mem[74] = 144'hf782fdc006af08e20a8bf078fd85f43af4c5;
mem[75] = 144'hfa6ef300fe9ffa4c0a3cf0bbf4910a20f60b;
mem[76] = 144'h0cfff7e5f9bdf504fe950b390975038df428;
mem[77] = 144'hfeb4f9f4fd8bf494f2bcf9f5f4cc0d00fe30;
mem[78] = 144'h0292f3f600a60707fc820b3dfafd02630852;
mem[79] = 144'hfee003defd9ef56903d60a50f1d502900d11;
mem[80] = 144'hfe6c0464fd4cfcbb0ba6f9d4f51d06d60987;
mem[81] = 144'hfb36f834f8eb04dffab908e4f0d601f3fe51;
mem[82] = 144'hf5cf0429051ef77bf681007ff743f197f4ef;
mem[83] = 144'h04f7f3e80d2e0e3bf26e0076f36efd38f8c9;
mem[84] = 144'h0035f0b609c2ffbe06fd0a0e00aafd36f851;
mem[85] = 144'hfa660673fff8fcb607b2f8a506fef1250e82;
mem[86] = 144'h0f3cf882f64cf4e80b25f830fa2005a1f49e;
mem[87] = 144'h05cf0ad30882f07df1faef9cf3edffa905a0;
mem[88] = 144'hf1930c14009e04be09d9f324fd1cf9f702de;
mem[89] = 144'hf63ff1470944ee4b069405690ca9f9c6fd8d;
mem[90] = 144'h0a8e0d1a0babf29bf46c0e4e02ee06870be0;
mem[91] = 144'hfe80f02dfecbfdb8f745fef0f49ff96502ff;
mem[92] = 144'h0135f6f804750747f1040b0c0d690b59f9a8;
mem[93] = 144'hfd6af4d4fda90e700326f14d004206b903a9;
mem[94] = 144'h0e75012e0e9f0914f8d50f84fcfe0f540632;
mem[95] = 144'h0c11fa7d0c5bfe2b09c50a26f5c30696fc85;
mem[96] = 144'h00740b160268055c08f7f37bfb81fe7c0f80;
mem[97] = 144'hf89008e308da086bf6710102fb5d0106f5a7;
mem[98] = 144'h0a7808ed0019f83f054dff82064dfa9cf7e9;
mem[99] = 144'hf8c6025609f3f2fe0a92f15909fcf1890184;
mem[100] = 144'hfaf30ca60a550dd405140059fafaf9d1f769;
mem[101] = 144'hfcfdf6f00d300913f4bcf0680d6b03e8f76e;
mem[102] = 144'h0f6ff8e5067e0653f843fa08f5fb0bf30d54;
mem[103] = 144'h084b03f5f1c4fb1bf3bcf2ed0abbfef3079c;
mem[104] = 144'hf1e100f5f5b301b60e2aff87eddcffe10a0c;
mem[105] = 144'hf3d701ecffdef280f4fc03190621f6a402e5;
mem[106] = 144'h0b4e094b0077f1280b4ef966075df6bf08ac;
mem[107] = 144'hf02b0636feb3ffff01390d2df57ef450088d;
mem[108] = 144'hefa6f639ef79fd89f337f89cf3f1f129f675;
mem[109] = 144'h034e0571f882ff65f965f83fff84fd3dfe23;
mem[110] = 144'hf83a0c62f5b1f5f4fa59f084ff110a1c0043;
mem[111] = 144'h0d85ff63f73bef4c04c20becf2b80b89f00a;
mem[112] = 144'hf7d607d80e9dfe040dc4093cf0d30d56fde1;
mem[113] = 144'hf2cbff9e0e9cfc9e08ae01b0f8d2fc2ef407;
mem[114] = 144'hfcd1078d0333f3fef5bf04db0f560756f288;
mem[115] = 144'hedfc088f073ff8230b4bef310108075c00b2;
mem[116] = 144'h0567f00bf5040ceff6f8fc64eea609ac0b5d;
mem[117] = 144'hee4efb42fdb70968f2af0497efa5f1bc0b2e;
mem[118] = 144'hf7da0d840c280f2df8350dcb0a00059c0790;
mem[119] = 144'h05ebf0a9edd8091e07630939ef87fac1fca2;
mem[120] = 144'h0065f7b60195ee830592f8fff38406ad0329;
mem[121] = 144'h04faf6e6f09109aef90f0a52f374026305d5;
mem[122] = 144'h0b8f057c0dd1fa6ff4c800540505f78205ed;
mem[123] = 144'h09baff940562fcfb00d4f8280907f895017c;
mem[124] = 144'h033cf5fdf8500c52ff4dfb99efb2fe320e9c;
mem[125] = 144'h09c509dff8e7f4a0070e0cb70057f1740930;
mem[126] = 144'hf032ff9d0114fca70886f4a30e36fd0efd64;
mem[127] = 144'hfb86f7ad0a690a20f43df78f0e3affedfef0;
mem[128] = 144'hf7630f3903b4f440f5c30f1306b00fa3fb06;
mem[129] = 144'h060dfa300602fcaef0c1f75f0414fd60f8ae;
mem[130] = 144'hfd7c0954f667f631fe5ef139f53bfff50b4d;
mem[131] = 144'hfa4407d90038f1a10ba30ea30a730763f68d;
mem[132] = 144'h03f1f3c609abf1a70cd8f47f04f30e710259;
mem[133] = 144'hf57009050bb0f296f20f093efbf2ffdffaa4;
mem[134] = 144'h002dfcfff246fc8bf8f0fa7606dcf0360dad;
mem[135] = 144'hfad009c5f8240092f8a9016b0818f48e00cf;
mem[136] = 144'h0b5a06d50bdf0f2b033d053a04840c67f4a1;
mem[137] = 144'hf68d0be90fd9f192f4fa0d94f2130419025a;
mem[138] = 144'h02030b3a069cf2c1fffbf05d0ba6fc4bffd9;
mem[139] = 144'h0e2bf7a7f75cf9880e9a099207d6fa9af56f;
mem[140] = 144'h0a41ffbffa34f655f9bf0d31ffc7f74207f6;
mem[141] = 144'h096ff814f9de0c8c05bbfd5ff285fada0610;
mem[142] = 144'h056ffbb50ad4f153f0ddfb240df2084af223;
mem[143] = 144'h04b1fc2ff1b7f2740fd6fe61fe8afe620557;
mem[144] = 144'h0cba08e4f4c5fe0c0da4f6f504390db5f182;
mem[145] = 144'h01950386ffc60622f13cf2d9f425f4330417;
mem[146] = 144'h010504c2f4650a820e0ef610042a017ef507;
mem[147] = 144'h073cefd101fc00e204fe068a05c6f400f103;
mem[148] = 144'hf717f90cfa3b0ce7f35706ee083cff8df683;
mem[149] = 144'hf2030657fd1a0e9108a00eb7ffbc032ef549;
mem[150] = 144'h0a78fcf10debf02006670ab0fa2bf8fa0a88;
mem[151] = 144'hf5e5f7d90cdc0a1e00a0f92bfd7df715f62f;
mem[152] = 144'hf7fdf49504630cccf78c0452f4a8f028fb33;
mem[153] = 144'h0ea00da5f48cefe0fb3e003cfb8d0c63f390;
mem[154] = 144'h07b907cbff3bffbc09820ab3f3a80a20f716;
mem[155] = 144'hf6da0056ffaff792f581f2920de3f91d093f;
mem[156] = 144'h0dec053309610ae9051d021e036308c80666;
mem[157] = 144'hf9130404f6b8f683f036f47af083fb210260;
mem[158] = 144'hfdecfc1d055d00200a19f76ff8d5ffe40d50;
mem[159] = 144'h04630483078d035a0dc4f7d10bad04680a50;
mem[160] = 144'h0d0a0df00ad30186f15c0691f591fec3f734;
mem[161] = 144'hf042f037f32bf79b00ed049cfbf7f95109cc;
mem[162] = 144'hfdc50d2ef0c207cd02900db80489f73003bb;
mem[163] = 144'hf701f60c02c4fdf1019f0c43f446038df758;
mem[164] = 144'h09920baaf42d001dfe81f8c1f56005380cf0;
mem[165] = 144'h04e2054b0c56f4cbf6a3f317f00df703fdc0;
mem[166] = 144'h0273fee803ff0424f0c90b080e440183f06a;
mem[167] = 144'hf329056bfc17f94803900c6d0bef058cffea;
mem[168] = 144'h0663f65500c0fefdf546021f0b5502a0ff10;
mem[169] = 144'h04580652faa5f553f1ca0898faaa0467fa77;
mem[170] = 144'hf0f30527fba50a530c6ffc6effde0a6b069c;
mem[171] = 144'hfee5fd650bddf8f6f453fa8d05c00094f273;
mem[172] = 144'hf0a60be8016408c5f2d4f9950fb6fad8f5d6;
mem[173] = 144'hf80701c7f830f85a0c9602a702ddf41af82a;
mem[174] = 144'hf4a60fa0013707b500c705d809e1fe6cfa02;
mem[175] = 144'h0f5ef0790449f32408c60233fa44072bf7cf;
mem[176] = 144'h034b07a3073cfca4f7b1f13ff1fb0cf40297;
mem[177] = 144'hfd49f1f7f92c0e5d0ddc0f3e0b94f0260559;
mem[178] = 144'hf01203640e1007ccf4ba02a5045df3ef00e9;
mem[179] = 144'h0e3efc16fd4df63afe3e0c4d050b09510f77;
mem[180] = 144'h0105f88808d0f60d009e0b3b0cabef7ff0fd;
mem[181] = 144'hfdb4fb6efba808a0f70c06160dd30e8c081a;
mem[182] = 144'h0047f9e3fa04f58feff7fe1102b103a4fa3c;
mem[183] = 144'h08dd0c51fb5c0abc0ae6faf50a70fc80f649;
mem[184] = 144'hfe95f50df6c20329f4b10672fd59f01701a8;
mem[185] = 144'hf6f10229f527f19207a7093601b8ff2200b3;
mem[186] = 144'hf27cfa8a043df709075800a50d86fceff3b5;
mem[187] = 144'hf1daf8fafe180a3009c0f7b3f2c409200bd9;
mem[188] = 144'h0455f60ffc65f1fe03420dacf9b5f09b0ba7;
mem[189] = 144'hf018f26a00def60dff59f258065ef66e0ad5;
mem[190] = 144'hff17f1e8f60800b00b60f54bfcd7f6750fdd;
mem[191] = 144'hf961f384f71bfdb802c3fb3300edf593f90b;
mem[192] = 144'hfb1af7f1f37afc9ff02b03b5fcfffc580335;
mem[193] = 144'hfdae0d3c011bf44502cef28cf6410d68f8f5;
mem[194] = 144'h053107900641f8660423f07e0f96ff86f61e;
mem[195] = 144'heef4fd1709d5f56df90d07b6fcdc08d7086a;
mem[196] = 144'hf1ebfeb50a7b03400244083ef95afd2d0005;
mem[197] = 144'h02ebf480f387fee80623f2eafd1607080c6a;
mem[198] = 144'hf0820b5f01d101eef2010d1efcde0098f919;
mem[199] = 144'hfe28f0d8045ffc9d0c77f798018ef330f661;
mem[200] = 144'hfbf2f6daf7e5f7d50746f5200d96f154f4a1;
mem[201] = 144'hf7ef01fa0bec04b80f280313f317f351f973;
mem[202] = 144'h01e1fef3042902be0d1ff3a2f67fff10f8a5;
mem[203] = 144'h0928047801d10d2af9aaf88bf2e8fa59010a;
mem[204] = 144'hfd2dfad8f6f3f64d08820bdcfe330af505f0;
mem[205] = 144'hf8ad01e1fc2f0615f438f69bffd4ff60fac0;
mem[206] = 144'h0a0cfeb6f433067a0636f7e10d69f0d10426;
mem[207] = 144'h0ae8f9810ea9ff64f8e6f0a905170f8e024d;
mem[208] = 144'h028b05fcf51607ec031a0193fb820283f801;
mem[209] = 144'h07930bb3f0140025026af506efcf01fff42c;
mem[210] = 144'hf75406c301bcf21ef487f8fbfc270bf6084e;
mem[211] = 144'h07980ac0f368f14df162feaa0b64fa1def8f;
mem[212] = 144'h0866f40807750a3aec8ff734f37efc4e01e6;
mem[213] = 144'hfdd7fbdcfc7e057e0424f63b0d5df9daff44;
mem[214] = 144'hee890071f2700074f8b3f40df5dfef1ff352;
mem[215] = 144'hf6adf2d2efef07bdfc82fbee0c2c0304f191;
mem[216] = 144'hf5d0feb3f9c50262f559e4d5f9a5f8550742;
mem[217] = 144'hef73fde00a92f365033d05210d3bf1d3039d;
mem[218] = 144'hf920efb10c76f11af43e070a081cfe0bfe9a;
mem[219] = 144'hfe6ef0b4f0980889f5a8ff31081101d9f199;
mem[220] = 144'h021f004d01a2efcffd7cff29098e05fdfaf6;
mem[221] = 144'hfab000710944048e05afef460be105d6f884;
mem[222] = 144'hf686f6e6f3bc0742fc0a03bc0236f9dbfa27;
mem[223] = 144'hf305f77c0606089e00ebeed1f406f1edf127;
mem[224] = 144'h045a060ef97e00950c67ef9bf5f701cd04e6;
mem[225] = 144'h08e9094cf8f9f13603efef6f0de90b23f7be;
mem[226] = 144'h02ee0613f974f116f1def122f855048303ae;
mem[227] = 144'hf47d0cc6f2b3ef88f967fa080b3208dc0037;
mem[228] = 144'hebbe03fcf962fbbbecb509450153f1340952;
mem[229] = 144'hf1b30847fc120825f565fa52f5e6f829fb5f;
mem[230] = 144'h04cf0143f7d5fab40b39f013f570007d0b20;
mem[231] = 144'h0028031b04eef3c701b9efbc0795ef4efa84;
mem[232] = 144'he7abe60a07e2f518ec090011fc7ffcdcffa6;
mem[233] = 144'hf0dffbb40ae60736f6dcf996f212f1c20c73;
mem[234] = 144'hf963f7b4070df0c2faac09e2fe32f3a8f321;
mem[235] = 144'h0c84faf6020f0e490c85fc91eff701f4f6d1;
mem[236] = 144'hf17ef6eaef560f010963fd95fc80fc11f987;
mem[237] = 144'h0a5d0d0c0f12091a034eef300d3cfe28f72b;
mem[238] = 144'hf044053304630eedf1f1044f0e7af6ebf519;
mem[239] = 144'hfe5f05adf265f193f1adefaff2f503a80c8a;
mem[240] = 144'h0c5b088afd84ff9b021befd30bac0b0af1db;
mem[241] = 144'h02650d0602a1f9fa0d5d0aa90352fd4705c5;
mem[242] = 144'hfb710d6ff15df8c6f6b0093dfea5fe57f4dd;
mem[243] = 144'hf72502990006f52e09f1f7b30590f0caf7c6;
mem[244] = 144'h021e01e8f5890d59f2a8ff520d8709cc0ed7;
mem[245] = 144'hfd25f4750ee50da4fbb8ef88fadd0bf607d9;
mem[246] = 144'h0ab8f26afaf1063cf20b0a5fef78f01f0edf;
mem[247] = 144'hf88fff1cf8210b0004a6f92dfe1c0a35fd84;
mem[248] = 144'hffa8f62409a8f6fe050e0aa70aec007a0f15;
mem[249] = 144'hefd9fdaefb65fee2fa06f1f8fbae0c7b0e2a;
mem[250] = 144'hf76507a7faa80ddff41e0a4bf71a073df9fc;
mem[251] = 144'h09380ed3fa2df4d60dd7f31209def67804fe;
mem[252] = 144'hf69802800a870513f6380d8cfe8d0e34fa72;
mem[253] = 144'h097ef393fa16fdb00b0b073b0bd70dfcfafb;
mem[254] = 144'hf9780ad0f549083107aef5f5f60d0d7809bc;
mem[255] = 144'hf8aaf143068e01adf79507d0ff9a0dbf0411;
mem[256] = 144'hf2b3078900d8f2d3f4bff48202dcf8eb0e15;
mem[257] = 144'hf44d0581f54cfa46f6d8feeef75ffc8df1f8;
mem[258] = 144'h014b0ef20b5204c200af06b4f39bf462fe8c;
mem[259] = 144'hfd10067e00f70456f15cfde302f7f229ff4e;
mem[260] = 144'hf63ff3d7ff95009000def4e80854f00ff475;
mem[261] = 144'h0ee3ef3e0e5f028b01f70324f71cfba9f53d;
mem[262] = 144'h0afcfaf90b6cfad30cabfa9e0aa60a1f00ac;
mem[263] = 144'hf46c00b700a407e10badf4920afefdcb070f;
mem[264] = 144'h00ad03f101bcfb3dfcdd075a0b690c5a0f05;
mem[265] = 144'hf4870605f5e605cb0a240404efc50534063c;
mem[266] = 144'hf750f21e0ae9fe0dfe7d0364f25500cdff38;
mem[267] = 144'hf463f24fff4c0d5900300ca2fa69087df718;
mem[268] = 144'hf8e6f75b00c4f3b305f6f286fb780780f412;
mem[269] = 144'h0ef8fd64f83100690da601ee0055f285f523;
mem[270] = 144'h094601b504b201c40cc90818f93308ed0c39;
mem[271] = 144'hf3e9fe50fcbcf793fd92f102f1affd66fe7c;
mem[272] = 144'h013cfa30f8cdf80600130b97f0b80539f2f6;
mem[273] = 144'h02ef08d6f5700e580c50fefcfdf901adfff3;
mem[274] = 144'h08fbfa860318040c05520127fb75f48405d3;
mem[275] = 144'h02980c91f53b030ff475f03ef82709b8029d;
mem[276] = 144'h0cd20d66f8e10b030352f63bfe78010af016;
mem[277] = 144'hfc2609d9f9cef9b2ffcbfff6f062f05aff3b;
mem[278] = 144'h0828faa0f327015af495f3f7f8ea07fc01a2;
mem[279] = 144'h0459f3c1f0f3f9fe0410fe9dfa59f52efb06;
mem[280] = 144'h0f21f78ef04cf1e3049b0a1701a30e990e0c;
mem[281] = 144'h02aaf4fb0c2d018bf64a0a6ef66e013d01b5;
mem[282] = 144'hf4ce01e700720e83fc73fa220221076bf82f;
mem[283] = 144'hfa83fbe20ea9fd570043fd270be3fcf004be;
mem[284] = 144'h087dfc37ff2c061efb7f02050c46f8ed07e0;
mem[285] = 144'h0d1b00d903ce07d8f57e00e9ff5a0bff090c;
mem[286] = 144'hf7250852f24404b00e5803230895fc2602e1;
mem[287] = 144'h068bfe6a0e320c4cf82c01800cf8fcef003a;
mem[288] = 144'hfcce00260a65fe49014af7d10c400329faa8;
mem[289] = 144'h05aa04d50583f690f0db0b29061d02780f74;
mem[290] = 144'h01cff2f5f09601b2fdaf029309160f61f900;
mem[291] = 144'h0061fa49f32f0d20f7bbfc510435001ef01e;
mem[292] = 144'hf832eadbecd7071600b8e89af9a9eb26ef75;
mem[293] = 144'h0976f9e10c9b0ba30be1f894f08cf322004f;
mem[294] = 144'hf66f099c0749fe45041e0100fbaefe1800df;
mem[295] = 144'hfd710000ff3ceeb4fa830699ffea0510eb6a;
mem[296] = 144'h00feed62f96bfef8fe04ff6902b103fbf05c;
mem[297] = 144'hf214f60af531ed9df77dfbd2091a02bff08d;
mem[298] = 144'hf3370e5808fe092b06a60ebdff60f85bf5ca;
mem[299] = 144'hf1fa0b53f2a8fa5f0c3e0d4aefccf51af39b;
mem[300] = 144'hfa37fca7f91b05330035f5230c62f0710805;
mem[301] = 144'hf9dd045ef205f45ff8ebfac4f5ecf385f140;
mem[302] = 144'h0a8605c70e43f9f1f45ef1adf59df7dcf602;
mem[303] = 144'hfeb7ffabf51ff4c4f5ac0ec50002f558fe10;
mem[304] = 144'h022c086809590459f4b60096fdda04e104d4;
mem[305] = 144'hfd2ff5520215ff8308aefc0f0110ff580cc5;
mem[306] = 144'hf97009c90ddcf5b2f543f690f9bd0f1703fe;
mem[307] = 144'h0d70f571f0bd035b08ea0565056d0b8b0a89;
mem[308] = 144'hed19ed2ef29504560ae3f90c0c1e0365f2e7;
mem[309] = 144'hefd8f517091efa730a91ef91fa5a039a0abb;
mem[310] = 144'h0046f936f8d3efccf67af68406a00809fa32;
mem[311] = 144'hefcc0ab20521013ffc2ff9a50994f9b105b6;
mem[312] = 144'h0052f37903acf66007bd0a2efa91fc69fd17;
mem[313] = 144'hf166eebafc3ef786fae9f1fc0526f4cd0c63;
mem[314] = 144'h01120dd6fcf8fe4df22b024605eef8ba0421;
mem[315] = 144'hf24dfef70df401e0fe01fb91f7a5f951f36f;
mem[316] = 144'hfee4f682f0e20eb2023ff272f6490cf7feb9;
mem[317] = 144'h072302e105eef3cef12ff270f9e7f816fafd;
mem[318] = 144'hf7790226fd26fe830d9ff235f091f9d5f78a;
mem[319] = 144'hf713fc4bfd8ef001ee36fc6b059c0cb2f405;
mem[320] = 144'h013400bdf87b06aaf69e002ef09ef9540007;
mem[321] = 144'hf48bfbec0152fdf9efd0ffabfd650139020c;
mem[322] = 144'hfd4704caf04ffaadf484fcc206d0fdb40e22;
mem[323] = 144'hfbf9fec8fb14fcfbff6ffbaf04fbf429fd02;
mem[324] = 144'hf541feb9ed440c0fec7e03d5f7050000fc33;
mem[325] = 144'hf43f07710ce2f195035f04c1ffcf0079033a;
mem[326] = 144'hff00f8fbf38ef383f96604da0ad400f80111;
mem[327] = 144'hea02055efb3304e2f0e5eee5f3c2f15f0170;
mem[328] = 144'hf346f2e9efcfeafffb28fc5d088af124f31c;
mem[329] = 144'hff980bd6fac1f1e0022ff07d05060c250398;
mem[330] = 144'hffcafa4c0b630893f3a7057af048043d0f1b;
mem[331] = 144'h0ac0f1d508cff067fb85faba090308a20b77;
mem[332] = 144'h0bceff38077c0910f7eff271004b03e4096a;
mem[333] = 144'h0af30388ef640b8efd3efd81037806390913;
mem[334] = 144'h07b2f8e103c8f6adf07f0ed70d350c740118;
mem[335] = 144'h028e0454f144fe11f361f843f7d7ff8a08dc;
mem[336] = 144'hf6040e3f03a90fad05a5005bf2b1fa6400e5;
mem[337] = 144'hf77408370ebc0a39fd1e05a40168f393080e;
mem[338] = 144'h0d6af58b0481f8390b88006104a108260223;
mem[339] = 144'h02680cd8feb4fa71f8cc0169faaa08f8f4a9;
mem[340] = 144'h02baf46af6460537fafff300f85df9fc001b;
mem[341] = 144'h04eaf28c0333fa4befc0f78ef59cf6d1f5b5;
mem[342] = 144'h02e108e00a98053aff20fc3dfc32f93bf576;
mem[343] = 144'h051a0a32eccbf83800e2ffb2080aef79054d;
mem[344] = 144'h06c1066805a302d3f369f64deee6eeb50b8c;
mem[345] = 144'h09f3f74cf8d201eff7bdf22dff68010e0837;
mem[346] = 144'h0780f4ce05e6f5e408810e2205ff0b2d0a7b;
mem[347] = 144'hf9630ed2fcbefd910128035bf5150bfff9c5;
mem[348] = 144'h0353fecef034f19b0d380c4405e7fc8c010a;
mem[349] = 144'hf84708fa025f0394f15105edf643efd80b47;
mem[350] = 144'hf117f638f59af7ddf056fa32efda0b110c42;
mem[351] = 144'hf19d06390971f8bc0026fbecfa66f374f5c8;
mem[352] = 144'hf2dbf579f33f0dd4017ff8ea0ed5f604fc21;
mem[353] = 144'h0e7befa8041cf08f02faf26df58e085107e5;
mem[354] = 144'h0c54ff64093c0a99f8ab0a170acb01df062e;
mem[355] = 144'h027ef5ffef64f035086e0233f093f1510eb6;
mem[356] = 144'h0396e9080039f73f09cbfb98fade063f0727;
mem[357] = 144'hf862f75afb4dfda0f7980bcb011ffbeb0d45;
mem[358] = 144'h000203170874fcc9f017fd4f06b8fba00113;
mem[359] = 144'hf4afecbbead1f6c1f007fc0aff580652ed1e;
mem[360] = 144'he1a6ec4e00be0c07e935fbc9eecc00410012;
mem[361] = 144'hfb56f545f33f0112ee0afda60245ff500c7e;
mem[362] = 144'hf517f2ddffc30e06ef28ffee023eff750337;
mem[363] = 144'hf611fb22f187fbbcf6fbf81906510b8f0f6b;
mem[364] = 144'hf1bdf7adff200ef3fd1bf1d809c2f06e0d2d;
mem[365] = 144'h088eff4e06d60faa087009aa029ff104ff0c;
mem[366] = 144'hf6c3f94c03380ec3fc3102bafe6cfceb0378;
mem[367] = 144'h047ff3cbfac60c0c0bc90a650247f3bf09ef;
mem[368] = 144'hf0410d050570f2f3f48cfd2f0bb2f3320897;
mem[369] = 144'hff3c01aafa58093bf64b004409bd04b10636;
mem[370] = 144'h0c240e0f00d9083cf7f9051900a808360f50;
mem[371] = 144'h031e0f0cf834f6ea0bf40efa05e802a80cc6;
mem[372] = 144'h01010a850726067bfd24f50cfd84f463f369;
mem[373] = 144'hfd42098cfcc90640f560099c0c08f53902c0;
mem[374] = 144'hf9c0f301086bf701f14d067f0c1cf52ff76f;
mem[375] = 144'h05aa068403090a44038ff03cf220080ff0cb;
mem[376] = 144'hfd7afe8df2f30d45f16009190c5b037af318;
mem[377] = 144'h007b0a8df787050e08ed0a4ef9eef351f4cb;
mem[378] = 144'hf47b09e6076af96f0c97fd0401fef5bdf672;
mem[379] = 144'h046afc9af5910d29f086fd38f2740d8c0f2c;
mem[380] = 144'h022cfd8bfed701fff6c9039df46af2c5fc0b;
mem[381] = 144'hff8df4aa0ca1fa6af113ff1bfe3ff9d9ffc1;
mem[382] = 144'hf8abfd84029b0d5206b108cefd3d036df57d;
mem[383] = 144'hf75e03d0f0de0d4b05a3090ffd2f08f20d2d;
mem[384] = 144'hf1de0802fb160e82fc1afd330380f91af909;
mem[385] = 144'h0a43fdbf0099014c096bff6b09d4fb14058a;
mem[386] = 144'h0f0bf46af9510bb20cabff61fc340f3a0cc5;
mem[387] = 144'hfb4ffcf5faa5fe2401fdf848fbedf17d0392;
mem[388] = 144'h0beff92507b9f77df8f4f85dfe47f3f206bb;
mem[389] = 144'h00a1f926069d0c2af2d9fd610461081d047d;
mem[390] = 144'hf0ab0795f2e9f37b0beb0d2103e0fb92fe38;
mem[391] = 144'h0020f1c4f8a7fcf2fcf3f4c1061cf7eb0998;
mem[392] = 144'hfc21026201ecfa1c0aa405390abc0b10f7e5;
mem[393] = 144'h00a6f3f60dd3f13fefeff72efd3e0dad0cc6;
mem[394] = 144'hf31e057af2d30d4101cbf03e0f7407e4f86c;
mem[395] = 144'h067d03d30d42f8b9fb92fa9a0a350982fcc8;
mem[396] = 144'hfddbf3bcff95fe8ef647fd40ff770a02fafe;
mem[397] = 144'hf2a80c8df640079cf6a9f0580678f79f0351;
mem[398] = 144'hf4fcf46bf0f8f29d04f409f9f5feff3bfe34;
mem[399] = 144'hf6e1f313fd2afc43fb180af8057ef9aef7fd;
mem[400] = 144'hf9a1f9010566f535fc860ee7f032fb5004b8;
mem[401] = 144'h0197f12b0b7bf174f658097eff02f9dcf8e9;
mem[402] = 144'h080c051a041bfd3ff28e0a9e03a5f15704c0;
mem[403] = 144'h0388f72ceedefa5cffa5f00107d5f650fa83;
mem[404] = 144'h045a02a1f0f00122f57ff8a0f0d602b1fe95;
mem[405] = 144'h06c6039502c8f29bf70300d5fcc10801f9cf;
mem[406] = 144'hf060fa2f0671fd66f0f703e10ebb0b3ef78d;
mem[407] = 144'h049c0480073005dafe1b0a53eeeaf66d04b2;
mem[408] = 144'hf51a0569f3bc0c3d02c6099af64bf8190b5b;
mem[409] = 144'h0abc04cbf9950aadf49f03f20e11f1a20832;
mem[410] = 144'h0d68fe67f447f992f3830e84f5a50131017c;
mem[411] = 144'hfd6000160413fbcaf13efed2fd6bfcea0eb6;
mem[412] = 144'h0eab045cff5bf59afab8f011ff86fde2f239;
mem[413] = 144'hfba70d1003940df1fc3bf62705b8ee87fb45;
mem[414] = 144'h06e5ffda0f55f2c3018ef8a5f77f0b020a94;
mem[415] = 144'h0d7a09d7f862f811f5eff42f0ab106e80d60;
mem[416] = 144'h057d03abf9700ef10100eefef75d00a10d7f;
mem[417] = 144'h06fffc200fa20060f45902120727f8460287;
mem[418] = 144'hefc9f634fd9d071c036dfb0c02a0fb3b0f74;
mem[419] = 144'hf74604c904d3f40d05990a4ff5f5f59d0c59;
mem[420] = 144'hecf7f355ef3bfa910492ffd7f7d50937fcda;
mem[421] = 144'hf3cf0299000809d80d330a8601b2fd08f887;
mem[422] = 144'hfe45f728fe39f95602a3fa2ef54ff0ec0b20;
mem[423] = 144'h039feadcec3c0476035feff10678fa6a084d;
mem[424] = 144'hfd230260fcb2f6a0e8daebd6ed170424f6be;
mem[425] = 144'h08fe0c1bed6000b0fb4c005d0cf1f196f54b;
mem[426] = 144'hee7001a105cc07300400fe60faaafd95f10a;
mem[427] = 144'h0b05fc01fbcf0d1609650120f9a0f99cf383;
mem[428] = 144'hf336000df85a09bc067c0dd6fbef054ff2c8;
mem[429] = 144'hff90fef8f0810857f4450ce3efb107680660;
mem[430] = 144'h00310121029c04720866064e02ef08f80ab4;
mem[431] = 144'h09850a4a0deff7ba08a0fbe10a4ef224fb8b;
mem[432] = 144'hfaadfebe05c0031af086fca8fe960fa1fa92;
mem[433] = 144'h0e6e0ace0ac1fe3d038ef3b9fccef4ba03c0;
mem[434] = 144'h0fb90408017bf231fa6bf8b3011fff40f53d;
mem[435] = 144'hfbd700e30b04f2befa790c160e49f8110c8a;
mem[436] = 144'hffb0f9ddf4f4043805e501a20b82f8b60299;
mem[437] = 144'h03e6f8bf09eef2a4fdda0d9c07faf284f0db;
mem[438] = 144'hf19af77bf2e9046efac806e503f40ea2f17f;
mem[439] = 144'h0135022507750ba0089e003bf0f5f131f00e;
mem[440] = 144'h0145067b070902860e2eff78f6ecfe470afe;
mem[441] = 144'hf1e7f0a10ed908f8f67c071800a50359ffe7;
mem[442] = 144'hf66f0cf506f9fb0006c7fa000451f2b20ef2;
mem[443] = 144'h0c8a0ee3fa15f24c09a5f9bd0aaffae1fa26;
mem[444] = 144'h05c70240fe78033c0e530478033e09e1f80c;
mem[445] = 144'h021e05b50faa049bf8d7f8b7fea5f3b70dfd;
mem[446] = 144'h0d9bfa47041209d1f636016902bcfc2505ec;
mem[447] = 144'h0f580df3ff97f4f4f3e6ff20f440f41efaed;
mem[448] = 144'h0360f2f8fc61f779011208a8f1f1f08b09f4;
mem[449] = 144'h03bb0348faddff950d9c027a05eefa2109a6;
mem[450] = 144'hfe2d03a8f61a0e12fa1f070b0723f5940050;
mem[451] = 144'h06fbfa7efb97eec00cc3fad00b480122f027;
mem[452] = 144'hf9d20c43fb120e49ee0dff08f2e701430cf1;
mem[453] = 144'h04d2f4fbf3e0f51df43dfed8f859021efc02;
mem[454] = 144'h0a340a7b0272f1980c2af4fc04e2efc4f54f;
mem[455] = 144'hf42df5f101ce0339042bf6b9f7f7084c03cd;
mem[456] = 144'hf2b9074bf9d1f4110646fab6f2b205d1f605;
mem[457] = 144'hf60bffa2f184ff450b93f47c0731f186037e;
mem[458] = 144'h038a0bfd0b89f607f10605bff37f0282f5f3;
mem[459] = 144'hf3b0f787f02cf2fb01480e6efd6fff400fc0;
mem[460] = 144'h08caf672fd00f99dffc00292ffddf844f934;
mem[461] = 144'h0e860a26f023fe60fe3604e0fa1608fa0b1e;
mem[462] = 144'hffd10d3df89c0ca8ff56f5ebfb94fa720b69;
mem[463] = 144'h08e8f230f10f0004f84c073305f40f45fb17;
mem[464] = 144'h0f980163fc87f2270db702cb014106120932;
mem[465] = 144'h0387079607f3050104bcf4e3f4500a56f076;
mem[466] = 144'h006dfe1707d205da0a5d0ef4fbb5fb610413;
mem[467] = 144'hff23fbb009b908d6f303f37ef90f053af23d;
mem[468] = 144'h0c3d0772f81e08ab0322f022ed18065cf97e;
mem[469] = 144'hf530f6f8f7c5ef9f06b70c1d00010dcd09b2;
mem[470] = 144'hfa4201f40a32f27004fef9e6f50cff7e0c88;
mem[471] = 144'hf86bf9fb02b201b5fefdfe7b0a0a0dedf273;
mem[472] = 144'h02caf164f7e80e42f18bee990b4807dc05a0;
mem[473] = 144'hfd2702daf712fa31ff15fa3efd32f605f650;
mem[474] = 144'hfcc0f308fa4eefeb008bf5dd067d04ebfefb;
mem[475] = 144'hfa64f5ee0a020531ff810189f2640af70523;
mem[476] = 144'hfb3efe4f04ea05f3f62f0632f0c6f8dffd39;
mem[477] = 144'hf532f7eb02e80a43036bfcd5feb50564fa46;
mem[478] = 144'h0b5ef799fa58fdf5f522f6b501d909f90402;
mem[479] = 144'h0140fa5a0086065af61602a8f70cf532fbbd;
mem[480] = 144'h04af0ef7f69ef996f36bf9e6fa600ceef3fa;
mem[481] = 144'h04810dc80dfe002bf6d1fc92002bf742f6ba;
mem[482] = 144'hf2d80516f6cff84a0199fc05f3e50c6e0999;
mem[483] = 144'h0335f6740f4cf8e408e3f4c307f50cf2f71e;
mem[484] = 144'h0d43f86c010206a309600815f63e0966f854;
mem[485] = 144'hff63f4e5fb98fc310ec007da07e2ffaa048a;
mem[486] = 144'hfd38f751f481093df862f4e2f452fbff08a5;
mem[487] = 144'h07aa0e08f40cf2d7efe00531ffd1077cf8d9;
mem[488] = 144'h00a2f3d7f1180f33065d0d9a0355ff6af4dc;
mem[489] = 144'hf4470779f0eb0ad2f16d039f0df4f1890614;
mem[490] = 144'h0e66f2d8fff50fd3f5e7f91a08f2089706a9;
mem[491] = 144'h0026f3ac004404d90588036df309f305fd12;
mem[492] = 144'h02f6f451f94e0383fa3f0e0001d001e1f705;
mem[493] = 144'hf57907c0f942027c088bf8cf0e6cfc88fcd6;
mem[494] = 144'h05e0f99dff38089a0cc9f60cf1e2fc3dfbb9;
mem[495] = 144'h0f1af2480c7d071af6fa0b20fba0068a006d;
mem[496] = 144'h013ffe26072f0a08076d0cd6fe670bb3f509;
mem[497] = 144'hf1fbfa64055f07bd0d3b01090560f2350f9b;
mem[498] = 144'h091ffe4ff334078a04a2f7a2fbbdf236fd5e;
mem[499] = 144'hfccb0afafdda06c3fa87f52f081504eefab2;
mem[500] = 144'h074f0bf70d720af50523f0cb013bf9affa6e;
mem[501] = 144'h0c57f856f349059000200f48f4ccff340fcd;
mem[502] = 144'hf016f8ba0bbc07b0fc96f627f48c05f7f44a;
mem[503] = 144'h01dbf64dfa27f0260912fa5502b60d7afb1c;
mem[504] = 144'h083cf86a014ff7b3096708a7f1bd0209f250;
mem[505] = 144'hfe0502d602620ebd0e23fe0806a80b4ef407;
mem[506] = 144'hf915f8cd054cfd4ff65cfa67f05a0a5bfcd6;
mem[507] = 144'h0c99041805340a770ed1f0a10f6b0207f6c1;
mem[508] = 144'hf05cf3d2f60bf7b9f90a0ba5f24007090b5f;
mem[509] = 144'hf4fb0ef0f053f8e5f637f8b907bb03b3f5e3;
mem[510] = 144'hf70508ee089f018df8dafd71f09f093ff915;
mem[511] = 144'h0cd5fe5b0f990a020b3608f8010003b90673;
mem[512] = 144'hf75502d40a37f26c0efaf2f80230f3b9fd46;
mem[513] = 144'h0dcb07a3ff4c0e31fc130bf1f4abff920a05;
mem[514] = 144'h06ef0b3b0cafff440b0af7b309ecf2f6f1c1;
mem[515] = 144'hf5bff1bc0e3cfd5af287019e019603500a68;
mem[516] = 144'hf888f73cf6f9f7f9f9a003eaff19f0750b1d;
mem[517] = 144'h0f84f345073e08720deefc500c4e0f6c029d;
mem[518] = 144'hfce40c570edcfbe7f47f0adaf26a0175fb3e;
mem[519] = 144'hf12efdba048e00270863f4de047ef270fa5f;
mem[520] = 144'h01c0f592f65c06fff9ad0d7704dff77e0223;
mem[521] = 144'h0d970c6af9f1f16af966ff1a00cf099cf103;
mem[522] = 144'h0bf30057f2b604be062005c009beffd1f823;
mem[523] = 144'hefd50eab0f79f4b5056a0cf30343f7d40e7b;
mem[524] = 144'hf8890846f491025fef89fa8600dbf07ff8b0;
mem[525] = 144'hf97205d508cf08eb0b2d0d7ff2160733fd66;
mem[526] = 144'h0639f3e40b150715f204fd1af0cf019d0ce2;
mem[527] = 144'hf32d0481f55af4e8f2f6f66604ac0407f90d;
mem[528] = 144'h0582f2210d75faf001a3f921f0cf0e2905ed;
mem[529] = 144'h0b470b79f8e6096fefa8028eeee1f38403f0;
mem[530] = 144'h00bb06900a500b5d018cefc80c6af6910099;
mem[531] = 144'hfe6bfae0fc7af80aff240a29f2d7fc3def51;
mem[532] = 144'hf03a049bfe56fbf107de05bc028cfa6702b3;
mem[533] = 144'h0509fe2af828feb20a69f2b502f50385fcfe;
mem[534] = 144'h05a5ffa7f2260e3d05e0f4fa0c330c1500b3;
mem[535] = 144'hfbacf068efd40246ff170192071c09ed0804;
mem[536] = 144'he93ce5bc0cd9ea45f5ddf71eeb7605c7f813;
mem[537] = 144'hf7440cc1027502b5fe20f5360ee30751feba;
mem[538] = 144'hef57f9b7081b0643f73a07180d36f99cf7ba;
mem[539] = 144'h0e4d017a0d52068703df0389f870f39c0099;
mem[540] = 144'h0717fbaeef0d0c0dfbe8fa340092f65ef5b4;
mem[541] = 144'hf9060672fab1f36bee61f8eeff1703f0f927;
mem[542] = 144'h00aa01e10da7fba30359f9d5f29c0144071e;
mem[543] = 144'hfee8f043fee8fa1d042df74df8e9f06f0b53;
mem[544] = 144'h0b8df64c005bf40c057b0b26f16dfe0b04f5;
mem[545] = 144'h04e0fcc402bffdc1f66a07d8f9cafb95058a;
mem[546] = 144'h07c5fdb40c3ff972fa270e4afb1303aaf44e;
mem[547] = 144'hfcd8f13bf557f6f70372ef81f00cf9f0f736;
mem[548] = 144'h04c70b12f52dfa7aff29fabf01d8f2f1f4ca;
mem[549] = 144'hf34503e601a40030fed50a8a0bd8fcb0f076;
mem[550] = 144'hfc02084ffbce02c0f04bf5660a87006df3ef;
mem[551] = 144'hfaef062707b00a8cee270921f43904f00410;
mem[552] = 144'hfafb0a38f00b0045f10407adf356fd460c18;
mem[553] = 144'hf22f00a803bbfb65fd250bd2f53dfa580285;
mem[554] = 144'h0a9703b60998065109e102effec00761f9bd;
mem[555] = 144'hf922f8f3f63af35bfd03fca3f15df25e0d69;
mem[556] = 144'h03c9fed00d7a06580bd301470b18ff610afb;
mem[557] = 144'h091e058bf089fb8cf04af174f689f4eb01ab;
mem[558] = 144'h068a0c2f07c70edbfb9bfd6503520098f650;
mem[559] = 144'h00b7074604680ade0de703fbff7109ba09c1;
mem[560] = 144'h0a4af405f5def4c1f65503fbf8510bb805ad;
mem[561] = 144'hf945ff95fa84f26a0b4ff225fd62f0db09a8;
mem[562] = 144'h04f4039cf2d0ffa7f4ee09a6f066f8bbfbbe;
mem[563] = 144'hf19d0b68f4d6f6c700f800410897fc9f05e2;
mem[564] = 144'h06cffaf1f3a8019efacafc98fecfff99ff07;
mem[565] = 144'h029dfc6a0a88fd37f8760e8d01f8eda4032d;
mem[566] = 144'hf6750bad0806faba0d800721fafd05490139;
mem[567] = 144'hf52a00ebfd1bff11f6fef2f9f7420152003e;
mem[568] = 144'h06edfbabfbc8fee3eb300047f9c7fc6ceead;
mem[569] = 144'hefef0bf60a4f01790c250822f969052f03dd;
mem[570] = 144'hf7130ad9fefff6c000aff30f0717f2e30e61;
mem[571] = 144'hfb080c27fa820b800403f1b0fc68059dfdbb;
mem[572] = 144'h0ee3f9aff2de0382f50509caf0a1f6e9fcfe;
mem[573] = 144'hf66e0a8ff2b8ef77f149f0abfc0af17d0553;
mem[574] = 144'hf5e90b420b41ff710aaf085ef767fc68f64c;
mem[575] = 144'h0265f880f4b80a39f9310863f88ef02dfb44;
mem[576] = 144'h02e9f1160341f1fbfe850500002d0b87f048;
mem[577] = 144'hfaa204aa0e980dde0b86004e07c506b6f8ce;
mem[578] = 144'h038c04840667f7c403df01f2f0e907ed064a;
mem[579] = 144'hfe07f06907d3f23807a8f70501ff0a2ff26b;
mem[580] = 144'hf880fcb3045af9b2f30d045404120d5ef050;
mem[581] = 144'hf995fed9f8900d8403df0a650383ffb7fcb2;
mem[582] = 144'h0b6905e8f9310838ffc70a52f2bcffe4fd4f;
mem[583] = 144'hf143ead30706fad6f4e8f32708d10a320600;
mem[584] = 144'h03f50ba8ef9c006af592f10ffcfd0cdb0c12;
mem[585] = 144'h01e60517f3ee01ba04edf9910291f76ef1b2;
mem[586] = 144'h0201effdfb4bf47ef5be04adf962f6620292;
mem[587] = 144'h0179f9dcfa6401e50d32f840f5400beff29c;
mem[588] = 144'hfef1fb94f9acf61c005ef4c80041fcef0217;
mem[589] = 144'h0d81f774f1aefe4006e4f9710c5e092a0c71;
mem[590] = 144'h0225f5f2006df4f408440a3c08ac0974f486;
mem[591] = 144'hfa76fccfff85070d03db0c9e042a0bdf0457;
mem[592] = 144'h04b6f85bf64a066af15aff0c01e0fb44f408;
mem[593] = 144'hf238feaefddafc1902680c58f417fab404eb;
mem[594] = 144'hf2980c67f572f40ef857fc5a0b1df9c7f425;
mem[595] = 144'hfea9f6b10d8108eaf4bcf641f1e3fbed0acc;
mem[596] = 144'hf9c70e27f09603b4ff7d0829fe770b020db1;
mem[597] = 144'h02750dcb07370becf809f0b2fa4c055bf7c0;
mem[598] = 144'h0a89ff2c0bb1068604f0f9fefa01040dfbd1;
mem[599] = 144'hf9690d150ce5fc96fb3a05eafdb4f55defad;
mem[600] = 144'h004dff64084afee5f3b000c9f646fa31f9fd;
mem[601] = 144'h0e4ff00cef71f31f02a0ff2f083705d6f9b6;
mem[602] = 144'h04740eb10de9f762040afa44f16f0d73f577;
mem[603] = 144'hfa63fecc07f504ce0209f7b2fc0e0e9ef727;
mem[604] = 144'h0f1efbf5f6c2f26afa360399f2d40f220d29;
mem[605] = 144'h0ed0fccc0af90f4206f4fe5c04e500a0f73c;
mem[606] = 144'hffb105a304faf76e0b7bfbf7027ff60cfca6;
mem[607] = 144'h0ba20880f833f8530e150725ef66f397fbc6;
mem[608] = 144'h0d44f75bfd21f2c4fc4ff480f7b504300871;
mem[609] = 144'h00a2f5dd0ec7084801edf37b0cd7021ff0ef;
mem[610] = 144'hfc0e0fcb0aa8f79a0f3704e00e10087d0925;
mem[611] = 144'hf14bfb390b87f99308b00739f7d70c70f552;
mem[612] = 144'hfcaffc370f7b08e609f903fbf8def563f347;
mem[613] = 144'h07e4f646ff3d02a6fad3f6630c48f23f085e;
mem[614] = 144'hfa47fd28f4e40093014bfe18f228f6370268;
mem[615] = 144'hfb60f6b202e80abf0f6802c4f2f00f6eef7a;
mem[616] = 144'hf3d506a3f4def7650bf00dff0e1ffb250f6f;
mem[617] = 144'h0691f5770f4e072af0df091f0c0b0c0709e6;
mem[618] = 144'h0bf90b00f6af018efcc509660c2a00a7f182;
mem[619] = 144'h009cf2d8f64afdf6f48ef63afc990e080841;
mem[620] = 144'hf5e40745fb1c0263f767fc9c0eae0e5af557;
mem[621] = 144'hfd69fd79fac0f41608820126f311f46e0009;
mem[622] = 144'h0b8cf49af6c0f76c02a6f46ef78df271f2a3;
mem[623] = 144'h0d810d4a02850366f64f027ef89706edfe8c;
mem[624] = 144'hfd66fb1c0b4603b9fb610e2f0d140b9f0aeb;
mem[625] = 144'h031ff6c4055709b3efcd03c3f6b60486012d;
mem[626] = 144'hfcd0074e074cfb76f4f90f340866f817f19c;
mem[627] = 144'hf22e0b66fc4ef15f0836f53a0a1008f2fdb3;
mem[628] = 144'h01110d0b0c490c10038c0519f29c0c5df3ee;
mem[629] = 144'h0a9009fcfc65ffcc09190a1cf822f20b0b74;
mem[630] = 144'hfb62ff560e17f328fdad0910f277fecb0b13;
mem[631] = 144'h0140f566f505066f0b0aee06fb8fedc5ee4a;
mem[632] = 144'hf2aff1cd0d08fbb0fbc10d63fe5b0828f7ae;
mem[633] = 144'h0d36fd710c82fa9e0045f430fa44034e01bc;
mem[634] = 144'hfeaaf2bcf2e50dc9efb5fb2d0356f792fa30;
mem[635] = 144'hf9e10acef9cb0066f690f3dbf58aff89fdb2;
mem[636] = 144'h0913fe2cf672f9410694fc950a1306050cb9;
mem[637] = 144'hf188f50206d6f6520684fd7af0d2f7d6fd9b;
mem[638] = 144'h0cf30231f78306d6fd2ff09a0f4206ea06ea;
mem[639] = 144'hef9ffc9a0c7a0d5bfaf7fa69fa27f01a038f;
mem[640] = 144'hf93af43efdb9f58ff92d0c2e0a3ef08c07e6;
mem[641] = 144'h0715fced068b09baf403f274fbeb049800d2;
mem[642] = 144'h05ff002f08d405f8095406d70ede05760a18;
mem[643] = 144'hf9afff300e58fa800b02f2e8f1ea09d7f8d1;
mem[644] = 144'h05c3f25008f605a8f3cf08e80006f33e0641;
mem[645] = 144'hf185f9160a15fadcf754f9f7f2c803a4013f;
mem[646] = 144'hf74301e70158f355fc810d9a06e8f2f60aea;
mem[647] = 144'h044f07a6eefc0194031302c70b39fb6bf190;
mem[648] = 144'hfd79f0f9fb9ff67d059afcdffd1bf338f0dc;
mem[649] = 144'hfc9cf0bdfb01f9d400d60297077bfcf9f62d;
mem[650] = 144'hf5c20c2601eafce5fb2df89defbffd42faaf;
mem[651] = 144'hf51702dbf4b30563032f044afb2a02480329;
mem[652] = 144'hf684046809ae0be9fb8909e80518fea2f4fe;
mem[653] = 144'h0884f381fb09fd0bf0f20c330a9f0a740f2d;
mem[654] = 144'hf46c0014046605aef3ca08870a6bf2ab049d;
mem[655] = 144'hf231f13c09690817fb42f258f2d3f2fa0339;
mem[656] = 144'h02780e4c0d5904c20837fd2afd76f2410e30;
mem[657] = 144'hef2ff0290e67030df662fb28fbcc063e0bb5;
mem[658] = 144'hfc77f150086ef0f50c15f321ffaff4380bbd;
mem[659] = 144'h0e1ff59ffd6b0a58ff2efd6407e90a7c004e;
mem[660] = 144'h01b9f525eb6ff634fa10f68dff8aee44f547;
mem[661] = 144'h003401f4ff61f42cf2110a72f782fb26fb54;
mem[662] = 144'h0d5f09590a3af556f599fd6afc5a0dbd0853;
mem[663] = 144'hefc30d200aadfcf2f4a6f4e6ef73fe58082c;
mem[664] = 144'hef10030ffbabfe9bf91108e70497002e0a2b;
mem[665] = 144'hf1adf40c06d3ee1907e8f6e1f2dffdbb0c36;
mem[666] = 144'hf886ff07f4faf24dfa220b5c0e9bfcacfe0c;
mem[667] = 144'hfe51067b049ffb46f37ef534f936ffd9012b;
mem[668] = 144'h070802c3fb07fe9e0d390cf2f9f008fa0d10;
mem[669] = 144'hfae808c3f20208e3057d0d57fe36f2df03f1;
mem[670] = 144'h0bcaf3590309f3e4f3d1fcc6f3ec04f60820;
mem[671] = 144'hfdef03f4faebf8a4f328f9630c440a01f2bd;
mem[672] = 144'hf8fa005afbf0fff2fe6109ed0f1dfc0a0d6e;
mem[673] = 144'hf50607e30e07fa640a51063f0ee6f969f5ed;
mem[674] = 144'h0188f376f1d30603fed7fdb801c10e28f64c;
mem[675] = 144'h02f5f9480625f4ba02a6f51f0b7af9d70ea7;
mem[676] = 144'hfd89062e0d38f62e0e04f07f08cc04190538;
mem[677] = 144'hfc6ffefcfea804330b56f32c0070fcac0d61;
mem[678] = 144'hf4d900300a750669fa09f4bb005cfb89f4a0;
mem[679] = 144'hf3a7fe2502f1fd3d0afbf8350770fef8f661;
mem[680] = 144'h0a3cefdb0c010e97f7c800d6ff21fb610273;
mem[681] = 144'hf6fc04afee930152f418f2910e31ef1df314;
mem[682] = 144'hfd9d0d6c079cf8c706f50f01048af6e201a9;
mem[683] = 144'hf78df7cef6fd06500770f44df2d50e2906ff;
mem[684] = 144'hef9506580877fa34094b0643f17af049f710;
mem[685] = 144'hf13505f1ff8e0d9df3f1f86e0d48f5dcfeb3;
mem[686] = 144'h0843ff1d0cf2fa4f0cfcfd82fb52fcb4f644;
mem[687] = 144'hf19ef2fa073c00ebf73d00790c6702e4fdf4;
mem[688] = 144'h03e7fc690658f91a09cffa62027bf4c6f723;
mem[689] = 144'hfed3f1fb0aae07f2fc67f336f5aaf2bc0dce;
mem[690] = 144'h03c80b770383f85803a2062b04dffe3a036f;
mem[691] = 144'h082e0cc3ffb3f9e7f86bfbe5fbd6f203f4c1;
mem[692] = 144'hf5bf07c101c7fd22f278f31a0604f3fff32b;
mem[693] = 144'hfd35f1f30b8af4d1f0530e75f5c10142f2aa;
mem[694] = 144'h0411f68dfc85060404980995f8a40b6903b7;
mem[695] = 144'hf3b2f30af45e0b28f424f0740f31fef8f379;
mem[696] = 144'h0cc4fc53f807f4690a72fa90f3a4fe4cff5a;
mem[697] = 144'h0b3602fa0bc6faa8001100b6f723f1e4fa95;
mem[698] = 144'h0357f64d0e8ffabbf15d0ed3ffa1045c0ba7;
mem[699] = 144'h095b019af7acf7180050ff5701e4f139013d;
mem[700] = 144'hf7fb0b19fbeafc98f04d03ebff9401c1ffd5;
mem[701] = 144'h0138f32b0711f93e091a07ecf37a02660b9a;
mem[702] = 144'hf68f04a80d55ff06f380fb2bf052f8faf876;
mem[703] = 144'h0a79fdcffbb3018b003002e80e5ff8320964;
mem[704] = 144'hf175f7fe02d60a930949fbbdf77ff1150050;
mem[705] = 144'hfb93fdcdf4f7ff3ffa2d09d30c3704440f3d;
mem[706] = 144'hfd5b0d4f0cc00b69fd21faa60f23fb740fe4;
mem[707] = 144'hf853efe3fb7c00fcffaef581091cf8420ba1;
mem[708] = 144'h0e6bf4eaf8f6088bfde70104061af67601a0;
mem[709] = 144'hfbddff4ef405f40209cef736011ef216fb64;
mem[710] = 144'hf470ff8af8650b200722f74807170f44f596;
mem[711] = 144'hf7d1f15502e803d8f73401bcf4bcfd52f32b;
mem[712] = 144'h042dfeef02e1f3150b610ed509c2feebfc68;
mem[713] = 144'h0343ffef06fff70907b8060ef815f343ef52;
mem[714] = 144'h02780704f72f020a0d390711f5b5f8d6f746;
mem[715] = 144'h0ea1fb3cf5290d4efbe8f1d8f5aaf5a90854;
mem[716] = 144'hfd52f3a7fd0e04990b1102b3f6dc0b460ad7;
mem[717] = 144'h0071ff6ff5fdf8feff84f6b1028b08d1ff5d;
mem[718] = 144'hf00bf9ecfea7f660f6490c95036100f9f20e;
mem[719] = 144'h0e9cfc73015404d70733f29df5b4f085097c;
mem[720] = 144'h0fd3fbacf33a0a30f90b096f09ed09060935;
mem[721] = 144'h0e7301560a90007ff85f04540187f885fa99;
mem[722] = 144'h0b09057e008401790f030d7e0cebf56ff15b;
mem[723] = 144'h00aff53f037001360f6c0c1a09b1f2caff83;
mem[724] = 144'hf7d7fb53efdd092908cf0a87f56d04ddf39b;
mem[725] = 144'hf78103fbf3a1f31efe94f182f90501f7f0bf;
mem[726] = 144'hf4d8f0e5089e03b1f085f0d30baaf9c3fec7;
mem[727] = 144'hf042f6baf5f3f7b2f77ef2040bedf5c50791;
mem[728] = 144'h08e7f9170a2402f4f8b5fdf4f55df5970ea0;
mem[729] = 144'hf15c076b05d00ae3f17701e9070e05a50e31;
mem[730] = 144'h00310594f92303aa0da00207fc6706520140;
mem[731] = 144'hff270e530f4c081bf1710810f43f04d40eba;
mem[732] = 144'h09b70ee80662f817015d040f0dc8fcb9f9d3;
mem[733] = 144'hf6560fd0f921fd02f52b0024f83803330fc8;
mem[734] = 144'h0e48fa11fef20705ffbf016e0b390cb4014e;
mem[735] = 144'h0e5f0dd001eff934fdac037bf7a80bc1f831;
mem[736] = 144'hf691fcc2fd320e03f22ff323fe4efa6a00b4;
mem[737] = 144'h0d980361fed1ff5cf9790c7ffa000c6503de;
mem[738] = 144'h01a2feca0032feb904e0042ef0c4fff5f470;
mem[739] = 144'hf053084b04ca093bf3f3f65af54405200299;
mem[740] = 144'hfe2d047efd130313f4c70073f9b1f9b2f785;
mem[741] = 144'hffcafbe1f3cf09e4fc43028c0e730a41f12a;
mem[742] = 144'h0b51f0cb0a8c0902fafb075df55e0aa8f141;
mem[743] = 144'h0a41f90e0ceb0bdb04980457fa39f56ffc18;
mem[744] = 144'hf5a70ac7f354feb5fcc5f902fd91fae1f0c8;
mem[745] = 144'h0733f92c024606dbf8b8004f08bb0835ff27;
mem[746] = 144'hf7bb059cf7c30c7201a2010d0346f9ae00b7;
mem[747] = 144'hf559f33506c9f09a0e8ffedff645f5e40224;
mem[748] = 144'h0a52f63f0f380e64f231f57904c006d9f141;
mem[749] = 144'hf192f60c0b7209f00e4eff2bfc3df49506a3;
mem[750] = 144'h0801f49df578f0ad0f2dfdbffb9f076d00ff;
mem[751] = 144'h061e07170e86fbbffc700ac4040bf77e09c3;
mem[752] = 144'h036f0da40d97f002f1c10e74f7ff0a2803c1;
mem[753] = 144'h0ea8fdf5f98efd91fdb303e50ccbf99b00dd;
mem[754] = 144'h0a050ec3f82ef4e208af0dd40260fe78f722;
mem[755] = 144'h0a5af59ef6d8f1f1fa94015e06370e3cf01b;
mem[756] = 144'hf0fe040c0ffbf51f06290cfff5280011023d;
mem[757] = 144'h0f4bf86204e3f36cfd4a0cfbfb3bf97a047f;
mem[758] = 144'hf65102e2f89e0413fbe2fa79fcaaf1790b00;
mem[759] = 144'h074409f9f739f1d5f24a023d061e0b430408;
mem[760] = 144'h0592fe9201230d070a02fc5400380aa2fc16;
mem[761] = 144'h027bfb06053efc2bfe4df9d7f1f3f6390f4b;
mem[762] = 144'h0114f130ff76f58bfdb100bf04dd08e7f5ca;
mem[763] = 144'h0641f3d5fc76fc1bf1690617f05df2d3fc9a;
mem[764] = 144'hf465f18a05d4094d07090f50fc55f06103b2;
mem[765] = 144'hf89002a80a6eff7d023501420e73f8f3fa92;
mem[766] = 144'h0cd509e2f59df79df8cffcbc0e8a0c40f945;
mem[767] = 144'h07b0057ef4340962f9b7fddc024a0f080e99;
mem[768] = 144'hfb13ffd5f1c7047e0465effe0e69f58e01dc;
mem[769] = 144'hf659f27b00b9f5a1f626fd38014806cefea7;
mem[770] = 144'hfa17f28e0f17f82ffd3ffd7a0753f21e02a8;
mem[771] = 144'hf6a7ff8701470aecf038f4c5043b044bff0f;
mem[772] = 144'hf34d06290499f600fd92f1a506a3001eef7f;
mem[773] = 144'hfe0503010ecffafdf923095dfccd0416ff92;
mem[774] = 144'h0e4df67407caf3abf392f2b5fc890ba10101;
mem[775] = 144'hfbc50a6bf329fec5f3910bb5f0b8049ef0c5;
mem[776] = 144'h0668f64309e9054af0c80de0fefaf04b05e5;
mem[777] = 144'hfc4d05a00065fd930528fed00ebbf16a0076;
mem[778] = 144'h08b509e6f67809b00d1efc5d0b270a29f5f0;
mem[779] = 144'hf9c50003f28107cc0df8f9240b12fe26f340;
mem[780] = 144'hf93f0b900abff2970304fdc7f685f7c901af;
mem[781] = 144'h0cfdfca80c8efef60f58f4c506eaf7bf0532;
mem[782] = 144'hf088fbe00a95f1ac0876fc95fc0f0524008b;
mem[783] = 144'hf94ef44a05a8ff7bfdc400b7097f00ab0c45;
mem[784] = 144'h06c20364fc48f03afd7af92df47a05a00764;
mem[785] = 144'hf4f3f8fa0a8af8fa02100484feb4fa77fb5a;
mem[786] = 144'h0b73fc580298fc76f4a0f987f4d80c690579;
mem[787] = 144'h0439f8fb0e000d98099cfdb00ee2fcae06d7;
mem[788] = 144'hf1ad047900d70b4b09750a98014efdacfe4f;
mem[789] = 144'h0eb9fd07028207b8feb40d0c0a97f3f40176;
mem[790] = 144'hfb6103440394f726f54df7430073fa840d4d;
mem[791] = 144'hf3a2f3fa0d79fe03fea0f75cfab0fae20476;
mem[792] = 144'h07540a5a044ef004f21cf28c037304c2f67c;
mem[793] = 144'h0b57f0e6018cf2fff2da0ad2009801e503e9;
mem[794] = 144'h0155fa8cfa6ef2360ef6f4ccff3cfccf0fbb;
mem[795] = 144'hfaa1fba3f4580074f502f39d0343f98706f0;
mem[796] = 144'h0e90f211fea201380d53fd0bfc7906bff529;
mem[797] = 144'h0a9ef724f4eefaa8f1a70c9109760c1cf569;
mem[798] = 144'h00c40309f48f0548fd380994f591fd1d0a92;
mem[799] = 144'h05200bd303510da4f404f7dbf3f2fc5bf5da;
mem[800] = 144'hf0a8efdbf797f3630c60f044fdeb0b1cf1fb;
mem[801] = 144'h004df20501320c1103effdb20956fb75fa95;
mem[802] = 144'hf6e5f0720efc0ec0ff100bd2f13a0d020722;
mem[803] = 144'h02960b300b5a07e50657085dfa0bf65f006d;
mem[804] = 144'h0182ea4c04c8ff4efc2b0450fec5f57cf3bf;
mem[805] = 144'hef37f9e2fc6c0aa3f767f863f77208a5f690;
mem[806] = 144'hef53f2dffcdbf9a4fd2bf11cf534f97e06f2;
mem[807] = 144'hfd2af11c0721f924ee6e04a6093ff245046f;
mem[808] = 144'hfdf5e5e8fe6fef88ef5df20ffe2303bafc17;
mem[809] = 144'h0e73fbc708d2fffe0a290ac20bfe015df578;
mem[810] = 144'h073af0c1f4adf0a1f1200953ffed02960b35;
mem[811] = 144'hf578f2fe0731019b0fad064ef0b6ff2af4c9;
mem[812] = 144'h059df290f0fffca905a4058e0c13f6f3f4d8;
mem[813] = 144'hffb8fb270409032a08ebf7d5fbeeed4bff63;
mem[814] = 144'h0a8cf4780a3f06a106fef17bfe37fa180b5e;
mem[815] = 144'h0b12f11e001b077bf4350b59019c0989f351;
mem[816] = 144'hf2040299f744f366fd11fddf0f08082fffb8;
mem[817] = 144'h029b0710f82e0bee05aaf28bfb430290f274;
mem[818] = 144'hf39802ebf153006c0af9f08b011c09090024;
mem[819] = 144'hf34108ff0e5df35b0892fd650599f99e0e98;
mem[820] = 144'hf388f73df8e0feb807e00a6ef782ffc0f6b7;
mem[821] = 144'h00bef108ef9ff194f83a00bf0407093c04e5;
mem[822] = 144'h0ac4f74804d0f9b9f6600928fce10c2dfc5c;
mem[823] = 144'h0842ee370785077801e3f1fefc6cf5b6f47d;
mem[824] = 144'h048d0ab7047b083f0b26059fef9ff823fa84;
mem[825] = 144'h0f40fb9aee8001a0f2edf65fff490d5d0961;
mem[826] = 144'h0e01f254feba04bc05daefb0f03cf6fd0485;
mem[827] = 144'h0e2ff6f2f1d2f8bcf2dc0773f220fab0f822;
mem[828] = 144'h0846f5e400fef78ff0f3efd1fe2ef6180ae3;
mem[829] = 144'h078f0e73ff14f17c08720d4cff75fb18f2ca;
mem[830] = 144'h04d0090f05a6f25d0ad9f440f4eafc6e0db2;
mem[831] = 144'hf046f858fab901ca00a00aeaf5970c1bf85b;
mem[832] = 144'h0d5908c3fb6dfbbbf4dc08fb045ff750f758;
mem[833] = 144'h062bfadefb36ffa1fb1303eb0e860cc0fc5b;
mem[834] = 144'hf2be022df609f3d90596f4a6f143ff1a04a0;
mem[835] = 144'h074d0f4b03b1f3e6fc770b72f17105a9ff81;
mem[836] = 144'hf7a5fce804d5f019f80ff121f1fefb24ffa6;
mem[837] = 144'h0afcff870c5e01ad09e90443002a07a5036e;
mem[838] = 144'h0ab90a7bfe760d5ffb63fe1defdf00530374;
mem[839] = 144'hfa03f9adfaf209740ca5f241f23cf8b809fe;
mem[840] = 144'hf118fd490e7f0bd501ba06020e74054c0691;
mem[841] = 144'h09660678f8a0ffeafbf304730d4bf2a8f278;
mem[842] = 144'h0937039004f5f9b1f4d101ac0f61f7fb01da;
mem[843] = 144'hf703023b031204730a48fa110a05fbac065a;
mem[844] = 144'h01ef0a69f6e8fe4cefcafa9ef6aff6e70445;
mem[845] = 144'h0faa099103920a3d06caf54409e5f2ff009a;
mem[846] = 144'h0d9e04a2f92ff2950b5ef9d3f55a0a690b7d;
mem[847] = 144'h012405e3efe6f5f1f7e0fad9fac4f1df0e51;
mem[848] = 144'hf27104e60d83f7a901320cfe0350fb68fab8;
mem[849] = 144'hf9a00484f5a703630e920e380171f819f769;
mem[850] = 144'hf4abf06400a10d2efe0f0dfcfffd0975f129;
mem[851] = 144'hf998faeafc18f97109d703f2f12dfe87f0e3;
mem[852] = 144'hf79ef8f4fa96080f007ef9dc00f109bbff20;
mem[853] = 144'hf86703130e36fa2eff09f3fdf1570c3805c3;
mem[854] = 144'h00840c9f0796f1af05a7f1670cd9f79c031f;
mem[855] = 144'hfda103f8fd9b0c19fbab07f5fee80b49f35c;
mem[856] = 144'h058906c4f143f885f4bb04cdf5eaf2e5ef97;
mem[857] = 144'hff30fd6b05da0ceff9e1f708f9f6f68e04b2;
mem[858] = 144'hf78dfc8ef237048cf4c708a0f10202e4f305;
mem[859] = 144'h06f0ff7f0eae05d205a20aa905950bdc025e;
mem[860] = 144'h07d7f72607e4f589f43af892f6f6f037ff8d;
mem[861] = 144'h031703f9fff1fe76fb71efbf0a53f0cbf335;
mem[862] = 144'hfbdd07f10849f9bef8d201e802edfc6efc96;
mem[863] = 144'h0d1c0d8e004701edfec6fdf00523efc4f24f;
mem[864] = 144'hfa3500b40007faf10c78ff99fdb0fb5a019d;
mem[865] = 144'hfabffec6fb1106daf715fe6007e90dd8ff4e;
mem[866] = 144'h09a002c70480fe13ff4706b6f6aa0c03f634;
mem[867] = 144'hf582fe97fd09fb0704d9ff9ffeae0851f210;
mem[868] = 144'hed68eb9eef0eff9dfc4bf18aee54f6c2ee19;
mem[869] = 144'hf1070d4c0efdf3fc008f0874f784fd0f0250;
mem[870] = 144'hfdcff322f32905c608110e01fc990d370c3e;
mem[871] = 144'hfab9098d046cef29eb76f17df8f0091a0638;
mem[872] = 144'hf6c8fc690af20259e32df219f3c902ae0075;
mem[873] = 144'hf8caf965faacfd34f57702c4f51409a8f9c4;
mem[874] = 144'h0fae0e7bfb1efd10012befa7f5e200f10398;
mem[875] = 144'h0b2df8a30b51036b0e6dfd0bf1defbc40b9b;
mem[876] = 144'h0304eee4f37d056b03daf602041cffcf0534;
mem[877] = 144'hfe6af680efdefa3f0670f3a4091ef638f7dc;
mem[878] = 144'hf9320a0905200ae0fd3cfb8d0f74fe7bf4fc;
mem[879] = 144'hfc74fb9d00130023f132f0a003c206c00490;
mem[880] = 144'h008a0a17099cf7f3048709a60271f88307b3;
mem[881] = 144'hfa8efba6f5c1f46e07c402da057206ed0610;
mem[882] = 144'h0ec3fb86fae70c6cf4cdf9ceff37058207fc;
mem[883] = 144'h059d06e1ef4304740c20ff59fb39f959fe19;
mem[884] = 144'h0cc3f9270b81fda3f45c095407910a10fdde;
mem[885] = 144'h029f076c0cef09a20492fc79feb405d6fdbd;
mem[886] = 144'hf23af523f4c5ffa5fa4df96306e609310eae;
mem[887] = 144'h0499f008fb72edecfd10f0e2066af0720479;
mem[888] = 144'hf68df05bf9360ab2000ef2110e8aefb4f3c1;
mem[889] = 144'hfebc03920702066d034a0c7b0b710f43f914;
mem[890] = 144'hf9d50f3df6a601b1f64bfbbcfdb301f2f773;
mem[891] = 144'hf2ce0088ffd3fdacfee20b95f478f59dfac7;
mem[892] = 144'h0c8b088200beefef0ca90c5409f3fa6903f6;
mem[893] = 144'hf785fbd30de1f724f212f07c0bc8f6810c07;
mem[894] = 144'h09cd08c7f1e8018f01aaf743fc9604280e03;
mem[895] = 144'h0e88008afbb5f5290cf407200f0bfe08f1e9;
mem[896] = 144'hf7cf0eb6fb33fc62fc8a01df0cdefabdfd2f;
mem[897] = 144'hf402fa4d0ab602a3fc6802ddf675f014f45b;
mem[898] = 144'hf621f0d004bff945062c0a7704d2f23ff9dc;
mem[899] = 144'hf95dfbf3f9e60ae903adfc70fa80f1f8f479;
mem[900] = 144'hf59ef24bf1fd0f17f51bf2390504fbca08fe;
mem[901] = 144'hf5350b2ef4f90211f52c088d03fa051e0666;
mem[902] = 144'hfbd50d8101ba006ef05cf686f308f3190256;
mem[903] = 144'h074a04d8eddef3c708190d310af6f9a00cbd;
mem[904] = 144'h07a70b00022df4a2094100a8fd4703070821;
mem[905] = 144'hfdacf059f2be062c07b6ff61fe160495f433;
mem[906] = 144'h09abfa6a0c03fabb006504e8f78cf7100167;
mem[907] = 144'hf1410ac9f5dc0a2a091608d709c2f43b08ea;
mem[908] = 144'h0478f08ffbc9f495fafbffef0807037805e1;
mem[909] = 144'hf31a011efc94058b0443f584f284f78507d0;
mem[910] = 144'h0d31020d0e52025306d5069506af056a0eeb;
mem[911] = 144'h0e7bfcacfeb70829f5d3f336fbbcf6d60c99;
mem[912] = 144'h0146f9f2feacfd72f7ce07ecfbb9f2a4003b;
mem[913] = 144'hf2a8f32cfc3cf6350af6f7250aa20b220a6c;
mem[914] = 144'h08d50f49fb5f08d6f67209d2f18ef3fb07f8;
mem[915] = 144'hffd90d440834089b048309220df609cdfdf5;
mem[916] = 144'hfccaf34c06f1fb19f41b0b03ef0ef54903ab;
mem[917] = 144'hf92afdec01bd099dfc7bf5660ef6fc800ef4;
mem[918] = 144'h00990c5cfd2bfe57f4fe038df2930f70fac2;
mem[919] = 144'hf4fef4bbefbe01340caef69703fbf185fa8c;
mem[920] = 144'hfd48fcdef5c8fb6bf30ffb35f30bf702004f;
mem[921] = 144'h0d3ffab70e7e0ea2f7e7fd850b16fd740737;
mem[922] = 144'h075cf2a201abf859fae6fc59050bf6100bf0;
mem[923] = 144'h0d59fb1bfe9b027e081e032d08b7fea6f5ad;
mem[924] = 144'h0b840315ffb0040c0c370c0a00c4f9e808a4;
mem[925] = 144'hf9a502fffc160e1df4e2f9f204670ef8f505;
mem[926] = 144'h09520b770efcfb7bf89cf79ff917f6a8f89e;
mem[927] = 144'hf15201f50c9604def98009c9f9b805d20e9c;
mem[928] = 144'h088b09660e68046e0af3effaf73afe6ef41b;
mem[929] = 144'h0149fb8ef02ff1f9fbc505380b6905f80d94;
mem[930] = 144'hf0cff43a0b36f1b2057c0cda0b72fd9c0b43;
mem[931] = 144'hfca7fc8b03ea0624f004036505a7fc670324;
mem[932] = 144'hf000fa71080bf6140efbf537f5310592f561;
mem[933] = 144'hf6af01e4ff20f9f301fb0e7803a00c320000;
mem[934] = 144'h0ea50f23fa710a87f90d08c9089ef3490bda;
mem[935] = 144'hf84bf3b0fc6b05d4f201f42101d6024a0b6e;
mem[936] = 144'h0612069e0358058a0bc007e00e44fcf5029f;
mem[937] = 144'hf057fdd90035fde9fba40d8cf4800a73fb86;
mem[938] = 144'h06c6084a0c320c64ffaf01ca007d005f0a8a;
mem[939] = 144'h0cf204adf15afb5a0703fbf8f5b0fbf200da;
mem[940] = 144'h0c73f2250b0903de0e08f4b20bbc09ee043f;
mem[941] = 144'hf31dfd6102cdf2f4f9fd002f05fafc63f4e2;
mem[942] = 144'h04bd017af7a2030df3bb08f00146f7ef0e80;
mem[943] = 144'hff4e002cf991f180fb6503610cf40fbf0e2c;
mem[944] = 144'h00aff91cf43b09330e33ff40fd8cfe89f6d2;
mem[945] = 144'hfa28fbfef9c7f20b069df4eef14a01fb0a67;
mem[946] = 144'hf3a4019e015ef6c3f3f90491f143090bf32d;
mem[947] = 144'h0957f12cfe2bff450b76f59dfad5f811f386;
mem[948] = 144'h045b0740faa5ff26f77f0a2904ebf2560e68;
mem[949] = 144'h03eb03b00b840cadfc2b0b3308500b4a08c4;
mem[950] = 144'hfddd0606f6cafefbfd4105580d6300960e7e;
mem[951] = 144'h0e9906c70dbdf894fbdf0a60ff7af744f967;
mem[952] = 144'h0e06f14103cd047bfbde07150eb60f04f38c;
mem[953] = 144'hf066087f06d7fc430cf5f01cf1c1fba2074e;
mem[954] = 144'hf25bfccefb60034cff79f97806f4f7f8febb;
mem[955] = 144'h0c8307e00197f590f84e049607450a6efb43;
mem[956] = 144'hf5cff7ac0b5c0765f74bfcc9f8f5fc8ff2a6;
mem[957] = 144'hfee20a7c02f00639fd02f5260cb8034afb74;
mem[958] = 144'h00780be3f86605240dbe0476fa1e05af0e71;
mem[959] = 144'h046402890795f1f802d0f4bcf8e90d700bb4;
mem[960] = 144'h0d79f00bf220f89ffbbef7d7f8b5f0e8f952;
mem[961] = 144'h0f8cff5c0aa10e11fafc0877039afaaeff5d;
mem[962] = 144'hf5f60ba0058908c50305041e047f02da0320;
mem[963] = 144'h009ef4990d2efbe1f4f10f17f72602e0f237;
mem[964] = 144'hf3100b17ef7d0bfefaf2f572fe1ff3f70d6a;
mem[965] = 144'hf0d4f744fb6ef33d02e809f1f78ff6ba0ed8;
mem[966] = 144'h097906fa082206d2f907f68ff6e8f2a8072d;
mem[967] = 144'h05880e26f82dfc5902b7f73a0ad5fcdff0bb;
mem[968] = 144'h0a470d73f822f39df282f0caf9210b3902fc;
mem[969] = 144'hf57bf9ceff82f2fef16c053efaaef82a0bc3;
mem[970] = 144'h04f2efec0f58fcca0d67077af34e0327f462;
mem[971] = 144'hf315fac90d4e0aba055d0f0f0a9af962f7e5;
mem[972] = 144'h0c61fc45002704fd04720855033ff63cfb86;
mem[973] = 144'h05df006af064fc06f6630e4308e9fbea0ca1;
mem[974] = 144'h07d007e003f3f2a0014d0628fcba05250802;
mem[975] = 144'h0b0f0f73fdf8015f0a37f5edf73804ebf3b0;
mem[976] = 144'hf47cf2f506960af8f1e9f98efdcf0448fe65;
mem[977] = 144'h06f90903f8c8009e0bddf6aaf888fa7704ee;
mem[978] = 144'h0d8d05d7f835061f087bf35f0026ff1b070f;
mem[979] = 144'h0c7dfa990e60017df847ff3a074a01d0ef95;
mem[980] = 144'hfd260a38ef6f0197fe8004f1feb90c3b0bfe;
mem[981] = 144'hfd89f3680c750247efaafc02f581016d03ca;
mem[982] = 144'h0c010d4b0712fcc9fe8a0574fe28f2680d35;
mem[983] = 144'hfbcefb00f9a7030cf47ff214fabfff900319;
mem[984] = 144'hf95908ecfe6c060ef8370095041c0d7eff83;
mem[985] = 144'hff630ec001c8f0ac0c9c03cbfaf8f39c0264;
mem[986] = 144'hfd580a800a280e4bf14c0cacf5fef1dcfd51;
mem[987] = 144'h0bd60f1701e00f250dd0fd910dee0a670690;
mem[988] = 144'h0503094006fcf0da02d4f0fcfc15034704eb;
mem[989] = 144'h0d2bf9110213f25ef132003bfcb0f1c7f2a9;
mem[990] = 144'hf1720996f783093203dd037b008202f50902;
mem[991] = 144'hf0e60e7afc1602befeeef4b80aaf08210165;
mem[992] = 144'hfccffa6c0dca07acf58f0ddc03d5f1dcf7a3;
mem[993] = 144'h017e060308ebf4c507d7f4bf06a9f242fe79;
mem[994] = 144'h018af11df3e20d0402320d320273f1120230;
mem[995] = 144'hf2adf15bfef9028ff435ff820a390dc8f1cf;
mem[996] = 144'h0618f0ebf931f79ef80df386f9f8ff10fa2c;
mem[997] = 144'hf53af741031703f7fefff00cf59ffe9bf799;
mem[998] = 144'h097c06b90accf375f98ff266f56a01910544;
mem[999] = 144'hfa0e02f603c200a5022d0de1fee8f6ebf31b;
mem[1000] = 144'h09650d0407820bce0b65f701f38ff8eefb21;
mem[1001] = 144'hf1a1fb47f03ef9c2f0def7b5f17f0f46feca;
mem[1002] = 144'h078df9600b7cf8fd0b560e790e2a040f0586;
mem[1003] = 144'hf5de030dfffa05fcf2ac0badf6980e120876;
mem[1004] = 144'h04e105dd03230f3308330e2f00f9fba9f696;
mem[1005] = 144'h0cfdf60bf2aa09e70c060704f45300470f29;
mem[1006] = 144'hf23bff050897f54ff131f4d70319fbb2024d;
mem[1007] = 144'hf13bf90e06cc0680ffe60a96fe2b00c907e2;
mem[1008] = 144'hf8b6f998f3790a6c0208f64000cbf55ff86c;
mem[1009] = 144'h06e30b1b00fd049dfdb90720ff76fe99fd5b;
mem[1010] = 144'hf0e4fe12f14c036e057c03f50c1cf5c3f786;
mem[1011] = 144'h0bb70a0bfda7f171002806e0f915f107fc7c;
mem[1012] = 144'hf156091c0628f8670555efe0011a03820368;
mem[1013] = 144'hfb7ff62f07f1f119fff60295ff760d65029d;
mem[1014] = 144'hff7fff17f4d8fc4ff44e060cf3280d370ddd;
mem[1015] = 144'hf7d10276efeffde3fb7afd02f047ff52ec41;
mem[1016] = 144'h0c23fa8508cf0323f069fbbefc14fbdfef55;
mem[1017] = 144'hf6abef660ace0170077df8b7f7a3f9e4020c;
mem[1018] = 144'hf977fd1af56c0c690122f0ab0e2df454faf6;
mem[1019] = 144'h04c4f01006a700800223f313035ff0050309;
mem[1020] = 144'h03fe0726021af8a7fd040beafde7f64ef371;
mem[1021] = 144'hfedfffa1f9d90629fdc2f2df028003d00b2c;
mem[1022] = 144'hf8740fd1f48700310830f876f3cd0184f07f;
mem[1023] = 144'h0746f07602eafdf70d25fb0e0b69fad6f42a;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule