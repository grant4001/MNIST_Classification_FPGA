`timescale 1ns/1ns

module wt_mem7 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h09da0a5a0d2d09b6044ff5a9fcd8feea04d7;
mem[1] = 144'h012b01fdf7bff2c7fe8a072505e2f0cf007b;
mem[2] = 144'hf702ffb900f9f8a7f2a205a2f21ef4bb08c2;
mem[3] = 144'hf10a0136f3e6f0f3fdd70b6d00380734efc2;
mem[4] = 144'h0256ee5af41ff6ce0268fe950b310ae208b1;
mem[5] = 144'hffdff785f04f0aa503ad0751f852062bf720;
mem[6] = 144'h067f055600ae0e2aef92f1be012defe3fd9e;
mem[7] = 144'h06600c06f982091b079402ba0a85fd3804da;
mem[8] = 144'hf44cfd6e034e0258f430fbedfcb9f04b03ee;
mem[9] = 144'h00ea03bc0713fea1fc46efbafadcff54fd6a;
mem[10] = 144'hf611f9f7fe50011df658ffb3ef46f1620864;
mem[11] = 144'hf9a00ca5f44208aefd3502e9f09900070438;
mem[12] = 144'h07baf3940d2af43b03a002fd0c32f57cfdb9;
mem[13] = 144'h0a2ef50ff8f3fb6ffcb807f5001b021e005d;
mem[14] = 144'hfa2bfab40c8603c404cef6a8060cfe63f481;
mem[15] = 144'hf105fc58fee906c40c5701edf4b2f270f74b;
mem[16] = 144'hf42afd0af105f886fb9ef377faf2f8ec0ad2;
mem[17] = 144'h0a1aff6105dfff4a0142f02d07e4fcc9f715;
mem[18] = 144'hf3990783f684f6900298ff9b029801a507cd;
mem[19] = 144'h076c001b0203fad802ef03780c2801530ce0;
mem[20] = 144'hfeda071bf5a5061f02ecf9d20936fedd0397;
mem[21] = 144'h0bfffac90ce2f741fda7f23df4930107ffa2;
mem[22] = 144'h08edf5eafffafc770334f092f7fe0315ff03;
mem[23] = 144'h0eb5efd9ef59f339fe740a41098f057df452;
mem[24] = 144'h0d6bf554fa6d068d0c98f3dbf120f68000d2;
mem[25] = 144'h01d60b8e005d0774feb0ef63fe5ef7090aee;
mem[26] = 144'hf81e0fac084b0fd5f1e7f6660e360bd6091c;
mem[27] = 144'h07f1035404ea0cbefd6cf582f852ef640e5c;
mem[28] = 144'hf806fc430b4cfa7cf9db01daf17301330df6;
mem[29] = 144'h007c0145f7e2f06dff19f87d0941f8f3f4f7;
mem[30] = 144'hf90307460d75f505002df1c6f40e0121fe61;
mem[31] = 144'hfaec0684efa6f1d8082d0a42f229fee00e29;
mem[32] = 144'h0398f3e60bee0b64fbe2078b098903cffab4;
mem[33] = 144'hf9bc0c72f2b6f1e4f616feb7fc5f026ef6a5;
mem[34] = 144'hfbdcf36ef2adf30bf286fe82f11cefdeef67;
mem[35] = 144'hfe5ef29701800865fd24009af8fb0be501db;
mem[36] = 144'h0dbd0b0905e30e320c0101cd00e50f490d57;
mem[37] = 144'hfb1df98a0de4f619f9dc0248f5350670f890;
mem[38] = 144'hf0e4feedfcb4ef6aefd1f54f001f03edf8cb;
mem[39] = 144'hefdcf3ef0f20fcd0f031056ffcd501ea087c;
mem[40] = 144'h035df53f04fa082a0cd5079e0dcaedb0079a;
mem[41] = 144'h0b88fd06024b055fff850a50018d00b6feaa;
mem[42] = 144'hfb950a1a017606a200ce016f100708acf4ab;
mem[43] = 144'h0b2b07dd03d8fdeffeb6f7df05dc041efa0b;
mem[44] = 144'hff43f664f85bfa60fefbeebdfd3a0c55f816;
mem[45] = 144'hf618ff01fa45035ff243fd4e03350668ffa5;
mem[46] = 144'h056a0c52055ef5edf1e30abeff5603c90f36;
mem[47] = 144'hf708ef9efab50c5c03b0fd060ef70c61041e;
mem[48] = 144'h0a37efb5f8fc0019f01c035bf1370b2602f4;
mem[49] = 144'hf30af511020f06c0f51807530381f11cfea1;
mem[50] = 144'hf161f88f02320e8a04abf8730ed20367f1d8;
mem[51] = 144'hf13bf0e7f118f7f5fdc1025a0467ff3bfdbc;
mem[52] = 144'h0a760cbefc52003a02a8f8100a51f37a0bee;
mem[53] = 144'h0a72fa410d55055ef86f07c4057cef3a002b;
mem[54] = 144'hf1b2f54ef30301baf9af0509f19ef7540cf0;
mem[55] = 144'h0631f206f713fef0f2e4ff9ff009f0e90d63;
mem[56] = 144'h0ca30474ff7101a4fa4ffb320bb5fa8a043d;
mem[57] = 144'hffc6efd8fb7a022d0932fca307a70945045a;
mem[58] = 144'hf026fbd2efd8f295f2bd03cdfac401ff019f;
mem[59] = 144'hf252f6050039098303310328080f0c70f74e;
mem[60] = 144'hfc190c0a0a180f21011cf6db0a4cffa9f2c0;
mem[61] = 144'h03f009fbfe7a0d82f5900acb05380cd9027c;
mem[62] = 144'h09ac0e04f3830c68f306fb20f231f6e7f9cb;
mem[63] = 144'hf6e10b0cf82efb990759058bf351f40af58a;
mem[64] = 144'heef6f597f1c7f6b9f513f669f06df9e0fe96;
mem[65] = 144'h01a70613f770fc9e03f8feb8fe45f80bf0b4;
mem[66] = 144'hf959f4150700f87700d6082f0e770e0af219;
mem[67] = 144'h0386f8190f0bfc750a33055dfc6f0dc0fb0b;
mem[68] = 144'hf5d4f2830dd4f0bdf3470f06f40e03e0fa80;
mem[69] = 144'h0620f286f5bbf4a9f5120bf1fb9509aff77c;
mem[70] = 144'h040df3d8f1b10d220e300945f379f6b60263;
mem[71] = 144'hfdb90da7f066011ff55e0196f923009a0abe;
mem[72] = 144'h01740e15f6cb023df99ff7a0f6b5fccffee7;
mem[73] = 144'h047d017104480cb60b420d97f08909fd0117;
mem[74] = 144'h06abf9c1f8770669068608b404cbf4d7f545;
mem[75] = 144'hfb6cf1120e5af55b09c8f892fa6dfa550c66;
mem[76] = 144'hf91a08200d690d0b00b80012f58303da0525;
mem[77] = 144'hf5e9001201f3025bff92f40f09d507f7fef0;
mem[78] = 144'hf2e6f7d701ebf512064ff5dd0927f7f3f049;
mem[79] = 144'hfaa40abdfa61f7460986f243f8f3f9d1fd0e;
mem[80] = 144'hfc16f365f707f87e0c17f246f03efbbcf69a;
mem[81] = 144'h0bfd09a0fb7ffebe0d65f8c6f34305f4f0a8;
mem[82] = 144'h0c5af73b0706f17801cffba5fd5cffeaff9d;
mem[83] = 144'h0807fa940c7502cffa4af52309c10e51f8d8;
mem[84] = 144'hfeae0c7f0ba0f82d0874046bf6b6fc0c0a4d;
mem[85] = 144'hf6cf0a3d0bbb097ef00bf8e306c6f058045f;
mem[86] = 144'hffa6ff95fffff0d1f6a2f8f20ef6f626f23f;
mem[87] = 144'h0033ff63fa6d0580fdbb04a2f1c3f621fe12;
mem[88] = 144'hfa720296f934f79008a407c70121f971f6d0;
mem[89] = 144'hf90ff96ef023f4beff2a08dc04aa0d5001df;
mem[90] = 144'h08ac04b5fa5a09c805d5ff18f4edf1e1fbe1;
mem[91] = 144'hf66bf8d4ff28fa08eff5f9490ab4fa26f54e;
mem[92] = 144'hfe85f35df57af1870afaf1dff7d80a68f06c;
mem[93] = 144'h07ac0b7ef915f139f632f18d08060086023a;
mem[94] = 144'hf16600aff8490deefc4afb7102840df10c12;
mem[95] = 144'h081609ea062c0e8bf2210ab10381fe170a9f;
mem[96] = 144'h0d9ff727f71e0fa40de7f1030b75fdfd0849;
mem[97] = 144'hfa9efe2c0197f771f87e00a2fd37f18b0975;
mem[98] = 144'h0e0d0f2dfb260bb40c93f58300b2f9eef4c7;
mem[99] = 144'h063ef441f9be0b56fd2dfb67023af4930fab;
mem[100] = 144'h04b60e6406f50e9f062d0c520aa6fa1df58d;
mem[101] = 144'hf94d03c4f2f9f78d051a00f7fe28f9ff0791;
mem[102] = 144'hf21dff78f0b5038cf59cf4d5f6820cac0d56;
mem[103] = 144'h0e62ff17f99ffb54017ef5fd087ff2e60c76;
mem[104] = 144'h093efdd6f3ee0f730db2f4d7f58f0bf40490;
mem[105] = 144'hf91cfdddfc560fca0e8befe9fd9404fa0768;
mem[106] = 144'hfc72febcf0bc0219ff2bf09bfaae0767f096;
mem[107] = 144'h06f10239f745ff1303bdf000061b05d30489;
mem[108] = 144'h0a1afc06f92001e1fd4bf55c0e1ff55ef573;
mem[109] = 144'h0caefd860a6cf310f83d0d5ffbf2f1e90c14;
mem[110] = 144'hf5a2f6fb03f20f11fe28091e025ef5df0b42;
mem[111] = 144'h0eab0479fbe1fb90061c0bbe0d0bf878f26e;
mem[112] = 144'hf14c05f80de60ec3fb05f31ef8cff4bdf63a;
mem[113] = 144'hf8a8ff9409a4f2590f640ab6f822fad2f7d6;
mem[114] = 144'hf2fc05d7fb9d0de90e0b0c7200be019c0404;
mem[115] = 144'h06dff9a0097efea3fb220263f3d406cff4f9;
mem[116] = 144'h01710caef2c6fa900761013401d6ff94f068;
mem[117] = 144'hff09f73c0c28f3980491f40cfef704250cd6;
mem[118] = 144'h0927f77dfa9c064f0ef704dc079df166f74d;
mem[119] = 144'h0284fb9701caf01df19bfc0dfa61f4bb06a1;
mem[120] = 144'hfd480537f3c90bedf0990c380e4103c40bb8;
mem[121] = 144'hf27c03f1f53c06ec05bf0879091dfdbefc52;
mem[122] = 144'h0cfafe2004cafc6707a8f40bf822f9f9f828;
mem[123] = 144'hf3c2f442fe47fe7cfd3f0884f862f9780c5f;
mem[124] = 144'h0af400c907dc0a290dcbf16f04cc0ceb0fad;
mem[125] = 144'h0056f0d1f1b5064c0d5102f000c904dcfc7d;
mem[126] = 144'hfe5f07ab085408e509ebf5d9f75cfeecf39f;
mem[127] = 144'hfa61f040fe4dff1dfa140f9f005d0b140c83;
mem[128] = 144'h01f7f65d0a91fe59fc09026c0f38f27a07cd;
mem[129] = 144'h02b8f13ef8e8021e0bef05950dfcf20f0496;
mem[130] = 144'h0142f875ff7c004bf95af6280d7ef0d3fad7;
mem[131] = 144'hf979f0edf87af8c0f4650e62080a0859072e;
mem[132] = 144'h0c71ff69f5c300a306a2fabaffc6f6c30405;
mem[133] = 144'hf69505b003bc0fd9074efa41fce808eafb0a;
mem[134] = 144'h0300f803ff29fef7f20ff763029ff06e019b;
mem[135] = 144'hfb320767008005a5f907064f074b095ef2fc;
mem[136] = 144'h08a1faa4f229fbcef12d066af43a0eb00e52;
mem[137] = 144'hff2ef2350ee40a67f4260ba7f2a3f664f3af;
mem[138] = 144'hfe08f2540ddafb0e02d3f9a5f385f2b9f83e;
mem[139] = 144'h041603da02f10bb6fef40ebf04660b3bf1d5;
mem[140] = 144'hf80903360ef70399fb6709990f0607b8f5c3;
mem[141] = 144'hfd000812f956029bf1f5fd7a08560bfafc2d;
mem[142] = 144'hfe3605acfc020e9f01fef3c5f3dbf3b3fad7;
mem[143] = 144'h084109ae05270685f267f87508f5f047f9db;
mem[144] = 144'h099e0bb6ffb2fb090e20f2b2f5970411fba6;
mem[145] = 144'h0938fd07fc40f7a2f5abf8a3f577f0330f04;
mem[146] = 144'hf6ca08a90aab0ee40955ffaaf7a806daf7d1;
mem[147] = 144'hf3cdf7d90952085c0a9c0b7b0f8f06c90c5a;
mem[148] = 144'h0019f4da0a7400e302f2f128f297f0430ad1;
mem[149] = 144'h0af601380fd0f4faf78e04ecf17ef6170bb6;
mem[150] = 144'h0ddefb25f07bf0dc0238ff0700d00250030e;
mem[151] = 144'h0ecbf68cfd70f3540799f7e0066aff7a0b5b;
mem[152] = 144'hf7e9f099051df7dfff60fc8ef34cf49e0fb9;
mem[153] = 144'h057406840488f93c068f0777fd38f96ff89d;
mem[154] = 144'h044fff6af062fccc033c0672fdcf04c90930;
mem[155] = 144'hfd2bfe2af8b105c2f03c0912fe820fb2030f;
mem[156] = 144'hf0cb0bf4008ef526063cf443f6baf453f1c4;
mem[157] = 144'h09c5fdabfec2f6bdfadb0533f7010d6f06a4;
mem[158] = 144'hf0b808ef0660f80e0887fc36f323fdde0315;
mem[159] = 144'hf4b8fa46f8d3f06ff02ffdebf22efa0efcff;
mem[160] = 144'hfa7a07da0a81062cf6210dc20f6cf34ef394;
mem[161] = 144'h0d5d0406f56507a00a60f33d0b3d0c76f0d4;
mem[162] = 144'h0d44f6d0f942f1acfce9f1bdf3d4ffe305db;
mem[163] = 144'hf76df6760a3ffc53f007004b0daafb500dc3;
mem[164] = 144'hf19ffecef78901b2f2740a0ff00ef3bafc24;
mem[165] = 144'hf83ef0e4f7adf8c7f450f019fdcef628fc65;
mem[166] = 144'h05900872ff6909f804df063f01b7040a01ca;
mem[167] = 144'h0426f46cf56505720f810084fb8df24d0be0;
mem[168] = 144'h0e45f3ac051ef33a08c809c906baf922f4df;
mem[169] = 144'hf5a00696fdd006e8f68e09e3021b0b92eff0;
mem[170] = 144'hfd9702520cb2f9a7fe20036903c7fde80461;
mem[171] = 144'hfd41f263f344f05f02c6f48d04c9f4ebf132;
mem[172] = 144'hf6130a95f4450ca103ebfcfd0e410eaa0cda;
mem[173] = 144'h0145f914f810f481f26804de0f23059b0563;
mem[174] = 144'h0cc7f9eafae10497fca3f918fc140b4400b0;
mem[175] = 144'hfc970d6ff5b909270c9c08f2009bf9360e1b;
mem[176] = 144'hf89af86d0b290307fb0cf0d1f784fc47f254;
mem[177] = 144'h090cf848fdc30f90fcd7f9a8025b0ce4f570;
mem[178] = 144'h0bc5007cfca9f1c6004f051407a7f17ef5de;
mem[179] = 144'h0dea0c48f83b0eb006b6f0ba00e8fd1bfecb;
mem[180] = 144'h05a4fda1081bf21002c1f652f7a7fd69ff71;
mem[181] = 144'h04b2f707fd7600d400c10dec0dd1fce40846;
mem[182] = 144'h0ca40ecf022cf413f28bef190117f14d012d;
mem[183] = 144'hfe2c0654f755fe12f6a8fc4605f6f81a07c7;
mem[184] = 144'h062b0283f12cfbcbf356f2e5f816f30df399;
mem[185] = 144'h0015fbac0607f982fccffbe7063efcd5037b;
mem[186] = 144'hf4b2056907a4ff66f9bff9a1f61df51b08fb;
mem[187] = 144'hef78f319087106ca03930a91faf60f0003bf;
mem[188] = 144'h00a7f77504c20ea406ad0086f47002a00a18;
mem[189] = 144'h0b0106070a72fc85f825f01d0a9ffa9a0c26;
mem[190] = 144'hfbfc086df7e8056b0a5d059106a709e500b8;
mem[191] = 144'h0a7a0d3bfe58f608072ef7b2003efa6af2ff;
mem[192] = 144'hfbfff23c03290045097f00e7f02bf00f0cd7;
mem[193] = 144'hfd2d042a047bf51cfda8f75efc2b0b1af4e5;
mem[194] = 144'hf6580f88f6c408e10d78fd96fdcff1f80b47;
mem[195] = 144'h0464fbec0f4af0150be10d22f164fc89ff6a;
mem[196] = 144'h0ebcfebdff4301e0f1800d1cfc09098f0d4d;
mem[197] = 144'h0ad609e6f36ff5edf4a5f596fc1bf82cf6a1;
mem[198] = 144'hf3bdf27a05540d2af603fe71f41df348024b;
mem[199] = 144'h0f46f06007e205030782feae0efb02c9fbfb;
mem[200] = 144'hf2acf821f569fd1e09ddf37a048806f20790;
mem[201] = 144'h05a7f269f5390f980d9aff30096ff8e7f4a7;
mem[202] = 144'hf1ea06d0fee406900a84093b0cf70b45040c;
mem[203] = 144'hf325088f0064fe0d065604ca09f90222f89a;
mem[204] = 144'hfc6bf7270668f481f474f59005bb0f54f9fa;
mem[205] = 144'h071803f6f6c40d85f8a60ded0009f188fafe;
mem[206] = 144'h0a97f0bb02730677f3860578f1300d8e0222;
mem[207] = 144'h035f058909580c1c0498fd38fbb3f00c0253;
mem[208] = 144'h0c70080a0a55f894f74af716f6be03a2f222;
mem[209] = 144'h001cf53afc60f7a5fc4df8e1f8210a9bf518;
mem[210] = 144'h01080a990a4ff786faa0fa6c0c9af6b10430;
mem[211] = 144'h05b6041ffc82f907fbea012af98d050901fc;
mem[212] = 144'h00e4f121fc1a0721f1cbf9f00a25f0050d42;
mem[213] = 144'hfceef4ee073dfbc409110cb40af80856fa0c;
mem[214] = 144'h03390e6b07e0f1c40e2400e7049ef99b01d8;
mem[215] = 144'h0cc4052c0cdf06140bd10b470096068e066c;
mem[216] = 144'hf217fee9f97a0b740c5fff78019502340ec5;
mem[217] = 144'h0f7d0d900c7df9d5f21301030a9aff74f87f;
mem[218] = 144'h0183064a0692f52cf9770e5bf442f96009f3;
mem[219] = 144'hfb31ffc10afef96ffde1f85ff9700c8e0be0;
mem[220] = 144'h0bdff258f862fa1a0da401d4023ffc86feb3;
mem[221] = 144'hfe9a05d0085efddff73bf7ddf4d10d64f4a1;
mem[222] = 144'hefe305c2f679fb26fb5cf9c0ff4a02d90892;
mem[223] = 144'hf308f67dfece07590d01f760f96903640432;
mem[224] = 144'hfd60f6f40588f87bfd9bfd3301c9069ef9fa;
mem[225] = 144'h088c00ea0eb60dae0198f141fed7fd330d8d;
mem[226] = 144'h0c73f0d9f4660535ffed0cc7fc8ff0ea0b07;
mem[227] = 144'hfa9d0ddb0193f5fffba7fbe6fe03fca20616;
mem[228] = 144'h0338fca30208fbe00e9e06130254018e0e23;
mem[229] = 144'hf6530e9cf15b0e04036bfa4a0c2904970c8c;
mem[230] = 144'hfa12ffaf050b032206cbfb68f04504700dbb;
mem[231] = 144'h04d7fae2f628011ffde20e3bf800f9cd082b;
mem[232] = 144'hf9c60c07f93e06e80887f5f106aef73f03d2;
mem[233] = 144'h07f8fef9091102d5038e0bb70a4b09dbf63d;
mem[234] = 144'h0026f6120b54fb6afd71040708cc08790107;
mem[235] = 144'hf1a80c4af6070909f6d6f327fb5d0103f9fc;
mem[236] = 144'hf978f676f6380100f88df1bd076ffd45f8c5;
mem[237] = 144'hfdbcf52f0819fd11fd43f16908a80e8b04e8;
mem[238] = 144'hfe45f81b04cffbcef7b9f57b04f800eaf8f8;
mem[239] = 144'hfb0bfea501a0f7740622029ffb41f8ebf06c;
mem[240] = 144'hfab0044604650356f576fa0ef01bf0ebf764;
mem[241] = 144'h0bae007ff266fa16fdddf862f342fba70ddc;
mem[242] = 144'h0e170462047df2b3038ffe4f07c50738fc08;
mem[243] = 144'hf3eff392fec505c7fbe90492fce1015ef61e;
mem[244] = 144'h073d0c3702640ecef529fc0ef98e0b75f864;
mem[245] = 144'h0a8d0c0bfd1f0db4f11cf6b7f0c2092ff766;
mem[246] = 144'hfbe50c72fe2ef66ffffa0796fd1b09f3fcc8;
mem[247] = 144'hfb7ef2030d9bffeef7bb0387f7010141fec4;
mem[248] = 144'h0387f599f7c50b83fbe40a80f324f042f0a0;
mem[249] = 144'h09700e48fc79022d07c1f2f9f3b7017908e3;
mem[250] = 144'h04ccfdf4016ff7e3fabf0df20594f6730786;
mem[251] = 144'h0aebfea1f571f4d2f4cffe5d0fdb0aef005d;
mem[252] = 144'hfb86f16405da0345f4fd0c5a0ed80d25f549;
mem[253] = 144'h0491f4ddfd1ff9c40f350b1df5d106aaf8aa;
mem[254] = 144'hfd66023501f7f372f5a9f59af1e209e5ff6b;
mem[255] = 144'hf0ebf7f5f6eeff35fc46f8fff66ef51ff59a;
mem[256] = 144'h0273f57cf7a700350b6c02bbfe4309eafd87;
mem[257] = 144'h0492f64c07cb00f60701fbe4fa15f55e0f63;
mem[258] = 144'h02a3fc0cfedaf8250961f877efb10f1df0d4;
mem[259] = 144'hf0b20cd2f1d606e10e50fd3b09c70e250053;
mem[260] = 144'hf4effb850f41fb2f0a0ff806f17f0f7bf2de;
mem[261] = 144'hf645f4960cbdf29ef56e0433f51602630566;
mem[262] = 144'hf39cfc22f13a09a402dffb2b037b0a7702c6;
mem[263] = 144'hfe71f3f50bdd0a43fd640e01f4fe06500a21;
mem[264] = 144'h0bea0dd9059102a40bbd0e490326f4760b7f;
mem[265] = 144'h015304fa0cf6fc84f6abf9e70211f8a9f461;
mem[266] = 144'hfee001b90852fa910603f4070bdd045ffb14;
mem[267] = 144'hfac70c43f954fabbfba500af062dfeb4f12e;
mem[268] = 144'h03b2062af3bef792fac103c9ef75f826ffae;
mem[269] = 144'hfc5ffedf0da0f63df2cff09dfc16094bf26c;
mem[270] = 144'h0cd501faf2690b2f0482034208f602f7f20b;
mem[271] = 144'h04a700880e720d410f13f44208c1097afdef;
mem[272] = 144'h023a057505530e550dbff53ffe59efd5fed9;
mem[273] = 144'h0aa8020efdbaf56cf285f3d706c80e1bfdd1;
mem[274] = 144'h004afa31fe8e0db50f61f5e60e5103fafe1e;
mem[275] = 144'hf166f7d502b7fdcb038efd16035cffba07cf;
mem[276] = 144'hf737f4350e01f0c1ff230c9ef5c3ff4bf02c;
mem[277] = 144'hfa3dfea10847f4c6fbb60fb7f382f710f79a;
mem[278] = 144'hfdfd065ff1c50ddaf5c0f1c40f6c06b4f4ce;
mem[279] = 144'hf6c40033f098f05bfdd00e74f40c07e60b96;
mem[280] = 144'hf8b3f70400a40f5c0f5d08cdfd4608460265;
mem[281] = 144'h09bfff3e0b70f4ee0f0b0008000f08c2f9a2;
mem[282] = 144'hfe04f41a0947f0400bc201e0f637f7750dcc;
mem[283] = 144'hf6d1f2410093f7260101fbef0b2802110015;
mem[284] = 144'hf0d6f524091ff0610b91009ffa300819f152;
mem[285] = 144'hf82b01c2f14e032af6edfcc6fcfbf4010c65;
mem[286] = 144'h0989fb110518fae105b60450f54906be0b3d;
mem[287] = 144'hf6eefda4f98d041ff74704310524ff22efc8;
mem[288] = 144'hf6eafbc709bdf251f1dff067f0430e99fda5;
mem[289] = 144'h01f1fccd01fdeff2ffc6021e0c44f054048a;
mem[290] = 144'hfac0eea10bb60b3c0e22f82100600709ff89;
mem[291] = 144'hf0e8f0c1fa2ffb970ad70be302b0f7a0f8f6;
mem[292] = 144'hfc9806a60c2ef0f30013042909200fac0095;
mem[293] = 144'hfbff0a93024ef1f90ca6fb5100a1fd520713;
mem[294] = 144'h04e1f72d076eff65063b03f803f7f737f50e;
mem[295] = 144'hfe8209dcfe7b0c0bfd0cfab10d47f824f554;
mem[296] = 144'hf0e7f2cbfab2f94809f70bbbf730f4420b11;
mem[297] = 144'h017a0be9054705c1feee0d22098708760a90;
mem[298] = 144'hfd780c83ef58028604f1f593feecfd27fca9;
mem[299] = 144'hf2acf742f63f02fbf32af6dd0e8609befd32;
mem[300] = 144'h03b0f1ba0df50e0ff8c60ed7fdd3f71803b0;
mem[301] = 144'hef6c0bec004907fbfbfaf589f0e9fe4bfc21;
mem[302] = 144'h0d700afa091309b9f7a1fdd30e6ff0b5f8f4;
mem[303] = 144'hfd6af108ff44f385f9ff08f0f12af11ff130;
mem[304] = 144'hf31908dc0b13f88e0372feb80bd0fc50f7ab;
mem[305] = 144'hff8402fcf6530da3fe28feaf0774fd150127;
mem[306] = 144'hf7770374f4a90acf0bebfec3f203f6eff82a;
mem[307] = 144'h03610f36f3a8f7fef0d0f6e9ff8b086effc1;
mem[308] = 144'hf466082b0e40fb9a06b1fcf9f799fcfa0c1f;
mem[309] = 144'hf49cf3d2028ff910ff070ec0f35df70bf4e5;
mem[310] = 144'hf2380a40f42bffbefc8e038c0fa60184f9d6;
mem[311] = 144'h0bf102faf79a0e92fc9efdea045f05ccf4fa;
mem[312] = 144'hf965f845fe3a0636f1420b77f20ef49d0040;
mem[313] = 144'hff680715060d0cbaf597f28bf24e09450901;
mem[314] = 144'h04abf54e0805f3bcf507031cf06301d6fdf6;
mem[315] = 144'h02fa0b0bfd000625f8140ac602b3074c0777;
mem[316] = 144'hf9a504f8056ef1dcf7a2f6e3ff700d5f034e;
mem[317] = 144'h0d74f36dfacc0c340bbbf548f2c401e30e36;
mem[318] = 144'h09b5eff6f1b909dd0554f79d0393f101f23c;
mem[319] = 144'h0820f8cafd9efc8b04cdf7a9f7ae0769f40f;
mem[320] = 144'h0e5c0c900127f3cdf7b002aaff0600dcfcf2;
mem[321] = 144'hfa29089ef80803e90f4ff284f47501de0dc6;
mem[322] = 144'hf743f42ff91d0bddf8e1f604f41c0f11ffe6;
mem[323] = 144'hf39cfa48f0020bacfd66ffddf0240072fe4d;
mem[324] = 144'h02aff78df91d078f01da001c042b0bb80d3a;
mem[325] = 144'h0eadf540efa807a106960ec80ef006aff948;
mem[326] = 144'h0753f060fd5df024f0a0feb1fb360d5bf5e4;
mem[327] = 144'hfbeef99a070e023ffc39ffe2fb63f969f6fa;
mem[328] = 144'hf81902b20334fe36f7c5fa0a002ff3540905;
mem[329] = 144'h02beee31f3d5eeb0f7350e9c088c09d4f029;
mem[330] = 144'h04b909e8f4e2083600fe08b3f264f86c0a24;
mem[331] = 144'hf8c8068bfb3d05f3fef8fd9ff37807a4f85a;
mem[332] = 144'h0b3cefc4f9dcf278f166fd9e004a0903fe4d;
mem[333] = 144'hf23e0b620c440309fe73024aff24040af06e;
mem[334] = 144'hff95f7d6f09bf4360dd9fe430a89fb82f012;
mem[335] = 144'hf11b0ab40824f3f705ef0972f7180266f9a6;
mem[336] = 144'h0b44037006990776fb65f8cffa11ffddfa7b;
mem[337] = 144'h0728f98a08d30ce70d09073a0027f742f5bc;
mem[338] = 144'h00280624f086fd7ff386005a0601fe690d66;
mem[339] = 144'heffdf32dfa91fd19f9ad0978fb840dfa0eb4;
mem[340] = 144'h00b2fa1ef465f3610f7400d80a3e07540a46;
mem[341] = 144'h03ff06790a34ffecf0a603250a07f057ff28;
mem[342] = 144'hf736f449fe89f878072afc9af648fc52f76c;
mem[343] = 144'hfffafc76fff6fe1406030d8d04a4f65ff6d5;
mem[344] = 144'hf8580ec3f1e603e80b94f60ffb9a0169f0c1;
mem[345] = 144'hfde9f5680cf900e6efab031900fbfd5902c4;
mem[346] = 144'hf6a8fbff0ee1f25402080068fda90e10f094;
mem[347] = 144'hf9a5053e0524f9790ad00bca040c0961f79e;
mem[348] = 144'hf67c0dc9026ff645f06c0004f07b0d5a05fc;
mem[349] = 144'h013afee70f4309e2fa0eefec0b8df88f0df8;
mem[350] = 144'hfabbfcd8f49609880717fee6f643fd62fd98;
mem[351] = 144'hf27afd86f1fafaf0f9d0f62afc1d07980e6f;
mem[352] = 144'h084f040df50df024094e078d07d8033ef561;
mem[353] = 144'h08b201bdf522fc2cf3fd09e6f2f403f3f8ec;
mem[354] = 144'hef66fd5608b70205fef4fdc90e8cfcc7002e;
mem[355] = 144'h03f2fba005e1059ffc07f7280e51f1e90d3e;
mem[356] = 144'hf26703ba087d07410995094efb030b95fce3;
mem[357] = 144'hf9d40eb7fd4af6aef7edf2b9f17ff5d1fba0;
mem[358] = 144'hf96ff3590302f89903e9ff160bee052c00f4;
mem[359] = 144'hf72a0ef3037a0cc7fe6a0ac7fad60a1e082d;
mem[360] = 144'hf02909ecf83e051b0c6a05d0fadf0657f08b;
mem[361] = 144'hf87cfb2f079cfe3c0b25fe91f314ffbefa51;
mem[362] = 144'hf6e9efcd0c90f6c6fc6a0e03fec2018ff7ab;
mem[363] = 144'h093afac7f31ef7aaf1db071cfa3f04cf0a59;
mem[364] = 144'hf551f8acf18dfe17ee4a095d06ccffc7f888;
mem[365] = 144'hfc1cf647f5860d36f944fbac0f35f09405ca;
mem[366] = 144'hf1dd08450819f34c0af6f5dcf3b3016ff526;
mem[367] = 144'h0c4dfc0af1a0f487f9820555071bf4160aa5;
mem[368] = 144'h09920cb7f48bf957f23f069efc4a05d4f7ad;
mem[369] = 144'h04d40ed507bc0889f59cfc7ffdbff43d020b;
mem[370] = 144'hf529f3d80f6cf6a8f2750d69f46007ba0fb4;
mem[371] = 144'hfd6ef0c00ff3f57a0ab0006e017b081903f0;
mem[372] = 144'hfa22f9ee03e80c2609f7f9d8029104480e51;
mem[373] = 144'h0d4301df0dd30d85f30b06200d4907950922;
mem[374] = 144'hfe79f05efe7702e00fcd0c82fd9d0fa6fd88;
mem[375] = 144'h087efe4407e4fdbf0785f9c0fa10fb690956;
mem[376] = 144'h0aa4fe63f6160aaa0821f2b0010df1b70c0b;
mem[377] = 144'h0401070bfcb7095708b4fb9ff15c06960cf5;
mem[378] = 144'hfdd10b32fd5ef8b4f994fd61ff16018a0f6d;
mem[379] = 144'hf789f04d04d80c59077605dafb86f7440c00;
mem[380] = 144'h0f9a0535f167fc9bf983013ef416f5a9062c;
mem[381] = 144'hf8c2f4f6f77d0c780462fc49f246ff4cf95d;
mem[382] = 144'hf48ffb8a018e0abaf99f00abfd36f0c2022a;
mem[383] = 144'hf9f8f24f0d2bfee60a080eb80ae7fb3e0f49;
mem[384] = 144'h087a05330cf2fb7af7cefbef0c52f163f1a4;
mem[385] = 144'h02240e72feb90cc0f805fded03f4feb5f9bf;
mem[386] = 144'hff9bfdee01c0f9f70803f461f3c4fcec077e;
mem[387] = 144'h070cfee90067f4ce07600138f50c0396fb70;
mem[388] = 144'hf37f05b1fa1bf1fffccaf402f540f6fe0de6;
mem[389] = 144'hf11209200cda0a09f7d1f3cc0ec6fdd3f9b2;
mem[390] = 144'hfe40f7c5f24efa5b01160746ffd0f35707b9;
mem[391] = 144'h0580f4620c7508b10172f631078e08a2f849;
mem[392] = 144'hf82f0b2500b6fdf10a6a0dfdfd310a110439;
mem[393] = 144'hf3840d2601f1fc050e170a6df86b00ea07f7;
mem[394] = 144'h0868f061016f08a2fd9101370e5d04810a1f;
mem[395] = 144'hf3c2f0770e0f066afa050362fcef01abf4c5;
mem[396] = 144'h0b4c06a40cc3f44d08e606210a490e3ff8a3;
mem[397] = 144'hf6d3076df06c009a04c7faebfeaf069df40a;
mem[398] = 144'h01060df2f4f400baf3b7f13309f3fc740225;
mem[399] = 144'h0b42fdc903450891f101047ffcb908e5f568;
mem[400] = 144'h0a62fba904c408b10abd0253f1eefe0bfc02;
mem[401] = 144'hf0adfdb002fdfbff04a5ff6e0d58f7610566;
mem[402] = 144'hffbdf9f6fca8feef0db7f3b005f4f49b0e77;
mem[403] = 144'h0a8d0ff0f04e03770baf01e4f71e0275f3dd;
mem[404] = 144'h0c7af635f4a0068afaaff4470c9df5a903e4;
mem[405] = 144'hf973f6edfc9b04aff8d2fc980ebef0b20c6a;
mem[406] = 144'h0bb4023203af083702a1f7aaf6aeff0ef6a3;
mem[407] = 144'hfe1a04a6f65ff2450c7bff43fae5012a0146;
mem[408] = 144'hfdc5f93e0509ffc3027d0ddbf552ff59fef5;
mem[409] = 144'hf54900b70890fe5e0a19022a016b07c109e7;
mem[410] = 144'hfdbf0bd8f92700b6f51d08ea0e96fdda0ab0;
mem[411] = 144'h0d090721f0510c81fdb0f5c3f6980a91f3eb;
mem[412] = 144'h0bd9fecf030f059f03eef91dff8608280eef;
mem[413] = 144'hf17a0585effe0c5ff1580d76ffaa04eef528;
mem[414] = 144'h08990595fa36f82ffc6ef64004dd00a1fc27;
mem[415] = 144'h085efb68f6bdf3670c230e6500d9f6b8f388;
mem[416] = 144'hf47ffd5d05760554f566fa37042df48b0803;
mem[417] = 144'h0b980efbf70cfcd202edfe4bf02f0d83f390;
mem[418] = 144'hefdf00ea09b500e4ff5cf9280f3a03590032;
mem[419] = 144'h058af758f4430cb407450ad0f841013cf312;
mem[420] = 144'hfffefc4b056e007ff3f904580cadfd74f704;
mem[421] = 144'h0028fd62071b06710245f8be090104c20c5e;
mem[422] = 144'hfe8ff955f0ff0ddc09ca0ab3f6c7f1e20d42;
mem[423] = 144'hf0400b5afcd5f15500aefd2a0545fc0aff60;
mem[424] = 144'hf9d9f75309e30bbafe0b0d9deffffc840b56;
mem[425] = 144'hf87f0d41f48bf9420573f1490b9606e9fa86;
mem[426] = 144'h06fcf513f845fece01100d98ffba0b0505b8;
mem[427] = 144'hf0fcf842068b0712fa2c04a9f5950a88f89a;
mem[428] = 144'h0d77fb710097f335065808b1fde5f213f7ad;
mem[429] = 144'hf25ff4e90556fefdfefef5c504f102e1f230;
mem[430] = 144'h0d86feb80c9ff0f603a80d28fdc4f790093a;
mem[431] = 144'h0c4ff6d5f163fc7008f6fad0f152fcde06ba;
mem[432] = 144'hf8b90e6df325fa53035bf47e04370f790b1c;
mem[433] = 144'hfb6f0ddeff57f67e0454f6370fc0f6280a7e;
mem[434] = 144'hf51af2e6011cefd1fc3b06aefc9308a0fc2f;
mem[435] = 144'hf381f244f697065bf96605baf97ef8faf797;
mem[436] = 144'h0320feaa06aa06eef1f10a8403daf83f0dff;
mem[437] = 144'hf36e03e8fc9702c0059202d4fa99f3f1f9cb;
mem[438] = 144'hf7d9f6f50df7f149046108f4072a01a905c7;
mem[439] = 144'hf8f0031cf763f071f9ec0ac1025af43ff481;
mem[440] = 144'h05eb0b4af6caf89af5c2f42c07dcf20ef1a0;
mem[441] = 144'h04420d3dfcf701b00028015d0641f8c30538;
mem[442] = 144'h0737f6d20025f0320d93fc0ff04c05290b76;
mem[443] = 144'hfaf203c4efbb0df5fc02016ef8beeedcfe88;
mem[444] = 144'h0ad2fc4ef43d01e7f45efca7f5e8efee0784;
mem[445] = 144'hfe1f09330015fc6afaf2f7a3f746fcb2fbe4;
mem[446] = 144'hfa2dfa5e0b9e09d7f5eafe3d02f8fe98f8c0;
mem[447] = 144'heea0f6adfc070eb6f77903970886efe900ec;
mem[448] = 144'hf4af061ffb3afc20f7700142f2ebf166f6d4;
mem[449] = 144'h03b0f8a30e7dfcaff758f53ff72c0e99f66b;
mem[450] = 144'hfcd405ec0b4bfe0cf109f23009d6fb380a8b;
mem[451] = 144'hf74c0b8fff390f990dd8091dfaa4fd8501e5;
mem[452] = 144'hf910f1a7f41b00fe0e6af598fb65085bfddc;
mem[453] = 144'h0817f30df29a0400ffa5f912f844f45e0654;
mem[454] = 144'hf35a0410f977fd6a08bbf619f5f1f6aef89b;
mem[455] = 144'hf91ff194088c05a807edf78d080cf6dbffb7;
mem[456] = 144'hf0c6f294f6dcf8b404e100bb0dd4fc200098;
mem[457] = 144'hfa1a052f0a1c0637f1fef36d01500913f40d;
mem[458] = 144'hfd0d03450f8ef7eff70e0363fbfd0d670c9f;
mem[459] = 144'hfa520ed5fbfef1dc0e84fd53fc420cf8fb03;
mem[460] = 144'hf467f5aaf3b8fad90326fc50f5d501f50841;
mem[461] = 144'hf1430672f3aafd72fbd0efbcf375f5fef4ab;
mem[462] = 144'h0efb0f45f776f7e9f9fff05df18b0ce7f715;
mem[463] = 144'h0653ff600decf6970d2af68f0181033f087f;
mem[464] = 144'hf0cf0b73fdadf47c0e3c004aff9bfc8508bc;
mem[465] = 144'h03cd03c9fb8e0348f0e00c2809e008af0e5f;
mem[466] = 144'hfbab056a094e0d08fe67f9440c5bfdbafa1b;
mem[467] = 144'h01bdfd290ef7f5d3fef2f9cb0b570adff8a6;
mem[468] = 144'hf3c7f5e70620f5700963f318fe2afabbf99b;
mem[469] = 144'h0ee50c810db8fc5bf040064605b50eeff93b;
mem[470] = 144'hf0aa0bba0b51fe800a86fda5f9aefb95fdd2;
mem[471] = 144'h0e2ef2530fb9ff9b06fe0bba0b470c6cf94a;
mem[472] = 144'hf0fa070603d50b820ef5f1960385fdc6faa2;
mem[473] = 144'h0337ff620f1d02640592fced0b55fb5bf50f;
mem[474] = 144'h0a5bfb170c3cfed8fceffaddef78061affa0;
mem[475] = 144'hf36d0a12fac807e4f6700302f4a80c2a0a42;
mem[476] = 144'hf673026df4c601ce0b74f2940596efd10c2d;
mem[477] = 144'hf3b905cdfc8f0c5d00bdf4e903b10b54fdd2;
mem[478] = 144'h0f01098ef1b0050ffb14faab01a5f8fefddc;
mem[479] = 144'h064ffc6df211fb9af844f738081d0ee8f0ef;
mem[480] = 144'h079e0893f056f932052ffff6f0d10375fcae;
mem[481] = 144'hfffbfdfdf658ffedf75af40ff88a0b1cf30f;
mem[482] = 144'h057209d101ab0021028407e8ff1cf55df2a2;
mem[483] = 144'h0077099a046dfc38fb7c026901120f2df178;
mem[484] = 144'h04b4f384f10bfa4b0af0f5a0f12b09f1f09a;
mem[485] = 144'hf162fe57f728072cf75cf7030e930a5c0306;
mem[486] = 144'h016ff0ae073cfd58f096f9b80aed0c4af48d;
mem[487] = 144'h095ef850f0ec0031f0ae08a9f560f003fd42;
mem[488] = 144'h04d80714f2580cd90691f2cc05640a29f202;
mem[489] = 144'h0547f4e5017efda3fd1ffb38f1e400d20703;
mem[490] = 144'h06acfaee067509f70183f7f70a3ef4cbfb4b;
mem[491] = 144'hfe44ff0df017062003bff73bfd420c5ffd41;
mem[492] = 144'hf85cf844fe25f2830e2af247055201800bbe;
mem[493] = 144'hf16ff100072c0f28f84ef87af25708a6f344;
mem[494] = 144'h07d305f2f2890a780ada0759fce900ecf201;
mem[495] = 144'h0899f504f523f9d40cd70d5df48c0ae5049c;
mem[496] = 144'hff39f83c0b73f4a9f95cfd33f6e7fa650981;
mem[497] = 144'hfa65fea2f7f7fe470538fc50f53ef4510cef;
mem[498] = 144'h0dc7f2090e5501f3fceff0e2034f07e302f0;
mem[499] = 144'hfb2704710414f1f20917fd070d0afa42f51a;
mem[500] = 144'hfb1a0b8bf42c0f2005dfffc3f0e5f86df64f;
mem[501] = 144'h0a56f8e30638fa710bfbfbbeefdd0157087d;
mem[502] = 144'h0e5c0029fd1d0e47f94efd49f9e4f49ef115;
mem[503] = 144'hffbd040001b6f728fe9d0cbefc7c0768ffdb;
mem[504] = 144'hf008efecffeb0e4001c1f02df9cbf925f2af;
mem[505] = 144'hf5ed02eef44cee4d0a93fdb30f02008e044f;
mem[506] = 144'hf6950365ef1c0530f5fbefde01360194053c;
mem[507] = 144'h00f304b9ef280b3d0d8bef6bf884ef59fb53;
mem[508] = 144'h0109026305c5fec30b5d086afe14f0970931;
mem[509] = 144'hf19706e0f73c048409650d27f128040e0956;
mem[510] = 144'h05a0016ff55bfd06f26a0b77feba00320527;
mem[511] = 144'h0cb7f578097403180178f170ee5508ee0445;
mem[512] = 144'h0518f6df0eccf43c09d9fe50f753fd700ae6;
mem[513] = 144'hfb37008a080109090bc80349018cf7e1f73d;
mem[514] = 144'h037ff2a20897f5eef6c4f058fed608edfa6d;
mem[515] = 144'h0b940e0a04a3ff9f0898080d0a83fe400f34;
mem[516] = 144'hf4c3f1470563fff3fe980d52fc58f1b70475;
mem[517] = 144'hf53cfb2e00fcf74d0502f4a602590619f869;
mem[518] = 144'h0ed4f4c1f46306e7f410fa0708d5f5ea0e55;
mem[519] = 144'hf0caf86308f5071af61f0cc30946fbd3fa2b;
mem[520] = 144'h0872fadbf318089a07e603150f7cf20ff44e;
mem[521] = 144'h0939f162058a0e63f83ffc390212f504f33b;
mem[522] = 144'hf0e4f7450c95f105fc7cffb4ef09022ef9dc;
mem[523] = 144'hf0bff66bf26708fe0d280554fe24fb1bf457;
mem[524] = 144'h09bd0d8e04d10dea0c190bf40556ff6f0b5d;
mem[525] = 144'h01eff5f30ef3f9def998f68ef830fa0b07f6;
mem[526] = 144'hfff1f2bef1c5f023fc3d0788f450073af5ff;
mem[527] = 144'h061bef8802f0fa00f2bef301fd62090ef60c;
mem[528] = 144'h0b66f35109ea07cbf3d509f0f4ea0804f475;
mem[529] = 144'hfa9002d7fc47f0720afb0b480715f4fd0675;
mem[530] = 144'hf08cf99afefef756f2fb0372fd9ff17ff46b;
mem[531] = 144'hfd62058a09c4fcc9044d0df1f242fdf00304;
mem[532] = 144'hf6c9fe88086ff7f3034df5bf0f14ffe5f68f;
mem[533] = 144'hf4dafabc067efefefff206b1fddff0e9faf5;
mem[534] = 144'hf062f81b087d0d07087c019b0c710c2cf7f3;
mem[535] = 144'hf66cf3f8074c0d6804de0997ff310fe9fd94;
mem[536] = 144'hfefaf89cf5630cb9073cf1d9f8030822ff5d;
mem[537] = 144'hfc66f120f1fc0f500a03f3f9074cfa07f3b1;
mem[538] = 144'hf7fff11004950230f44505500ab1f798f92b;
mem[539] = 144'hfe86f4d207f80757fb0af33df770ffbaf1c0;
mem[540] = 144'hef0e04360b01f2a702f8f7f1f9b0f12ff416;
mem[541] = 144'h04ab087af4160ee60bda08550e52f2cf08ae;
mem[542] = 144'h08460d4109490eedfb04fe29fe20f796012f;
mem[543] = 144'hf9baf3a80e42fd1106020113f3dcf4c30b09;
mem[544] = 144'hf00bf290ff8d02ab00be0bdffd8ff4a5f4c4;
mem[545] = 144'h05a20309ffb7f6780944f73604830b8c059e;
mem[546] = 144'h0bfc04dc0a320292020dfd6ff0bdf8d9ff47;
mem[547] = 144'hf905fd95f6e006c1f4810edbf8a80dd804c9;
mem[548] = 144'hf23e07c6fc0c0ee20e4700e1059f0312f41b;
mem[549] = 144'h0fb90c88f940f915ff8402b80a18f83af400;
mem[550] = 144'hf7f1f261065b0127fecd0397f8ed0232f549;
mem[551] = 144'hf91ef5160042ff45f79ffefcf29ef4ab00cd;
mem[552] = 144'hfd040a4cf6220177f9abff050a1ff9a9f093;
mem[553] = 144'hfce6f87efb00f302f423f6d2f78cfffc04b8;
mem[554] = 144'h0a2003a50d2d08a4f4540a53fb1b0f310698;
mem[555] = 144'h0f34fc2e0e3bfae20edf0e1cfe9df32409f7;
mem[556] = 144'hf965f9080a98fd810a4a043f0aa3f76a00b3;
mem[557] = 144'hfb9e06ff083d09a80b1c08e5f0a20b4c05fc;
mem[558] = 144'hf1efefa8feb0f9d1f3f50b0f005ff577fc28;
mem[559] = 144'h0b340f27fb380f81f49cf2c7f5de034cf2a1;
mem[560] = 144'hf021f4c408b9f6e0f248ff62f47b01af0fe2;
mem[561] = 144'hfa1b09c40bd90e57f412f9330ef9f501fb78;
mem[562] = 144'hf9450000fa8d0dc6f5bff7940191019cfe00;
mem[563] = 144'hfd470698f9a2f506fe6af1b00bb90ce60199;
mem[564] = 144'h062a0f72f6eafcc2f40a0b29f47afb37f66b;
mem[565] = 144'h01dcfa7cf7bffc0dfe580d1ff29af709fcfc;
mem[566] = 144'hf22d060106e70ff3f42205fa04df0f5bf658;
mem[567] = 144'hf061f22900990a9e010007cbf5200b65f7e6;
mem[568] = 144'hfbe207930635f122ff56f50d07edf4c20677;
mem[569] = 144'hfb39f2fd08ccf9be0a29fe72f03ff16eff40;
mem[570] = 144'h08b1f4c205a10149f2a0f1860f0afbaff3d5;
mem[571] = 144'h00a2074408a9f331f55ff2f3f06c03d4fddd;
mem[572] = 144'hf54a048901e3ff830f77faa4f629f7fd0e9b;
mem[573] = 144'hf17bfe6a050e03aef7b2f4acf5bc0f98f905;
mem[574] = 144'hff45f27ffb67fa47fead085308b90eaef296;
mem[575] = 144'h062efc1ef6b0fe82fe46fa49fd9bf484f062;
mem[576] = 144'hf45802a6f15409a5fde50217f27f0b5f0801;
mem[577] = 144'h05860cac0f8302150ee802fe0b8200baf4e8;
mem[578] = 144'hffdffd4cfce0f4c5f5bb085807befed9fa52;
mem[579] = 144'h08b2043ef5cbf447022c03e80d7b0b4eff04;
mem[580] = 144'hff58f302f41ef7a205a504d1fa3700e6f479;
mem[581] = 144'hf75606070f7a07c40cf90061fba9f43ef3d3;
mem[582] = 144'h046af47ef5cef008f2e0fb17f2aafadbfab4;
mem[583] = 144'h034402a4f92b0ac8f082f5a5f3f3f9250e60;
mem[584] = 144'h04290b9704b7017b04960da802b002d2ff69;
mem[585] = 144'h0545fe9bf75aff0d03d9f6090d06f160f91d;
mem[586] = 144'h0c03f519f3d5f82d010ef2e10305f9b50e86;
mem[587] = 144'h0be901b5fced07e6063e0d15f2a9f3cdfcd0;
mem[588] = 144'hf7ef01860389f4580cd904c904230c4c0ee1;
mem[589] = 144'h044d0944057a03b50ad0f2600249feca017a;
mem[590] = 144'hfb00fa22fb150baa0c8cf484f339f69f0322;
mem[591] = 144'hf52604bd016a0ae40e9a00f8fa4df08bf2c3;
mem[592] = 144'h088e0c09facc050b07b501990701f94bf566;
mem[593] = 144'h0cf50b780a990b480751fe45f46406a50d96;
mem[594] = 144'hf4090a1a02eff6e0f02efd0ffe58f443f18a;
mem[595] = 144'h0d0507b80b63065b08d506dcf871026c01c3;
mem[596] = 144'hf046038b02650a2a0d57f260f02ef37a0dc6;
mem[597] = 144'h08b8f4ddf0820041f4e70aa900e9f6a3fd5f;
mem[598] = 144'hfeba031df97df1b0f62efecf0b480a540e57;
mem[599] = 144'h029e058c04b3f8870613f3a5040befeef836;
mem[600] = 144'hf5e60806f795efff05c3f084fbabfcb6fd17;
mem[601] = 144'hf6a3fe86f67201ad092506d1f88e06e50e7f;
mem[602] = 144'hfb0709140dcefecbf4050ae50f6a08980c65;
mem[603] = 144'hf3f2f9fa035def47f19a001ff4b10def01e2;
mem[604] = 144'hfaf90a04f32d00ecfbdb021ef32af5a4fb7d;
mem[605] = 144'hfdf601e7fadb0939fc040649f2e70aa40bc3;
mem[606] = 144'h0d820e930cd50df5ff95f89d04cef76efe32;
mem[607] = 144'h0ab70afc079dfd7f0557052ff32804f40de3;
mem[608] = 144'h0bc6f7e7f2040216f393fbfbf2220e9df4b3;
mem[609] = 144'h06450859f7330084f184ff1f0c4bf9420b81;
mem[610] = 144'hf0cefe40f13100500092f5c7feac006bf24a;
mem[611] = 144'hf98af3cff36ff9260e8f09890ea4f1c7f086;
mem[612] = 144'h08a1f23e03a1f4f4f216f6b50cc803dd09da;
mem[613] = 144'h01d604eef8c1f2cc010dffb2f60af6250df9;
mem[614] = 144'hfd78ff560735064f04ce02060b9d0491f72b;
mem[615] = 144'hf8bd02b603bcfd750afffd0dfcaf055dfc70;
mem[616] = 144'hf48e0e0c0dc6f26e08abf1d10f530e930a57;
mem[617] = 144'hf316fe48f7b5f5bfef0309370290ff1cf359;
mem[618] = 144'h04dd0b5504ac0e9504480a80fcfcf5a90070;
mem[619] = 144'h0b29fe09f3200a430e73f5ed01080f3bfda8;
mem[620] = 144'hfd08fcf9ff0afe860167008bf70b0490f256;
mem[621] = 144'hf51d05de0b1106aa0e700f69f6c70963076a;
mem[622] = 144'hfdfff01000070d64017c009def9b0402059c;
mem[623] = 144'hf68ffeaaf172f1fc01530ceaf86d0d8a02e7;
mem[624] = 144'h0b7cefe90a530630f3f0ffbe039d0e15fb2d;
mem[625] = 144'hf79e0b17f14ff9a60c60f7e301f7061dfce9;
mem[626] = 144'hf1d90b9a025dfd75fc99fde0fb5ff03d04f9;
mem[627] = 144'h0e86f2c7fe35085e0e01f731f38bfaa80106;
mem[628] = 144'hf422f293feecf8bef6020cbc0b84f4bf0988;
mem[629] = 144'h0f2402a306ed0fdcff7cfd74071e0c290530;
mem[630] = 144'hfedb084b003d029efe850cf9fad40cbcf7de;
mem[631] = 144'hfa2dffe40906f06ff68c007bf49b026c0a37;
mem[632] = 144'hfbe8f1f1003ef30ef5f4f2a306ebff7bfb21;
mem[633] = 144'h0c35ff28022303a6f09f02340eadfc880061;
mem[634] = 144'hf9390b7508990252088cf272f7b4fbc8f253;
mem[635] = 144'hfb82fea3fc1cf7f0f906f3d7f864ffccfb28;
mem[636] = 144'heee4fa4b026c023f0b360997f79f0cfefece;
mem[637] = 144'h011a0f6d0ab2096ff56b03f1fd2004e1f50c;
mem[638] = 144'hfa8602080704fafc0d66f04408b10f340065;
mem[639] = 144'hf0dafb17090deff00882f0e7f53002960a2f;
mem[640] = 144'hf35a0d20f147f812f3a7efd20e870c27fdef;
mem[641] = 144'hf7e40f380762fd65f74c0a0a0d7202230e91;
mem[642] = 144'h081df3bffe19075bfe98fb66f78d08c7fed1;
mem[643] = 144'hf2dc0613f87808dff9bdf20cf71df7830168;
mem[644] = 144'hfc9cf391fe08f13d0f41fb0509ba0446fb36;
mem[645] = 144'h0b7df18304f1f202092cf3c8f1b5f000f43b;
mem[646] = 144'h06ba092af15f0f74f862f5c003abfe980dfa;
mem[647] = 144'h0c78f139f5f1f5f10c13fd30f4760ea10c59;
mem[648] = 144'hfa8dfdcaf3a705470ce6fe3709daf62dfac0;
mem[649] = 144'hfcaffdd5fac105a7ff7f0b7bf49c0048f193;
mem[650] = 144'h0cea0c24f653fa82eff407b9f725062006db;
mem[651] = 144'hfe340442f7c5f32704f6fbc3f9b80926f3fe;
mem[652] = 144'hf342f0d906c4ff95f9d5fd5af405022400e6;
mem[653] = 144'hfb7ef64afe5206090231f0a601650573f22b;
mem[654] = 144'hf671f68709adff58f1230609ffd505440c14;
mem[655] = 144'hf61efb9606ba03800597f6d9037c0eb708ca;
mem[656] = 144'h0cf8f8070353f192fff7f02dfdeb07230cd3;
mem[657] = 144'h03a7f9f2f630f9ddf619f1e9fcadf7b40340;
mem[658] = 144'hf458056b0f1afd5c014c0efb0cee0dc60563;
mem[659] = 144'hf6c5fba5fd5f05e8035e06f0f84c0b22f911;
mem[660] = 144'hfa2af31df2d10351f4dcfe67f3540e7cf023;
mem[661] = 144'h087def84fa940d3c0e1c037f08d30d68fb75;
mem[662] = 144'h0225fd3a0ecefab20269f87b0c3d07860bac;
mem[663] = 144'hf707f6e508e600970990f6c1000302dcfe45;
mem[664] = 144'hf44dfd040dec0a27f374f2160cf3ff5afd01;
mem[665] = 144'hf2e704ef0454fb9df765f3aa040c05530892;
mem[666] = 144'h0c0df9f00645fb3ef6ab0571f48e0d410bf1;
mem[667] = 144'hf710ef4efd65fc72f03900490c4ef91e0026;
mem[668] = 144'h0cce09200dda03fbf935fa4d082ff95501ae;
mem[669] = 144'h0d23f1900de70f8a0da4fe5af1e600920b95;
mem[670] = 144'hfd9e091df23b0ce2fd6bf3ed056ffcf707de;
mem[671] = 144'hfeff0ddc0cb8f2da0c8d05c2f3fdfa150b49;
mem[672] = 144'hfb96f4760dbc00ce0140037c0241fde2f3d0;
mem[673] = 144'hf5d609b600bef1bdfe190ccffbb4f5fbfd78;
mem[674] = 144'hfcee0057f3caf876fdd303ec0bd202effbb3;
mem[675] = 144'hf7b80ca3fc8303ba0c88f2cb010d0a2609d7;
mem[676] = 144'hfd5f0e4c014ffd9703ff0f32038b082df26b;
mem[677] = 144'h09ae00280c8b0aa1f0f40b6d09860897f29b;
mem[678] = 144'h0563fa78013802d0f4a401f5fa73073cffea;
mem[679] = 144'hffe805c5028a097df5eb0becf5640983f7ae;
mem[680] = 144'hf62c00bd04500f1e07540db0f8dc0741f5a7;
mem[681] = 144'hfee00a65f7ea02d2f56cf283efeffce40291;
mem[682] = 144'h0432f4510781068a09830dc407a40366ffa9;
mem[683] = 144'h01b3fc630524f6ff01def80af5bdf647f6ed;
mem[684] = 144'hfdaff9a0fdd305cbfb720b55fa5bf1d20921;
mem[685] = 144'h054906ca0527f014024f0005f6820bcdf5ff;
mem[686] = 144'h03b6f171fff6f862f5c30ddc010bf7f90e2a;
mem[687] = 144'h0d37f40d0089faf3ffa1fa1ff143ef5d0d47;
mem[688] = 144'hfa78f35d01ec03aef1ad0223f6adf2c60a96;
mem[689] = 144'hfcf802530cc007f7f793f97d09e40a8af631;
mem[690] = 144'h0d7cf615f1d0fceef0f008c30a9ff7e40adc;
mem[691] = 144'hfbc00a6d09d8f7d4f2560597fc840fcd0c54;
mem[692] = 144'h0fd9051906fffd310636f925fc40fa3ff432;
mem[693] = 144'hfeb4fe2a09520bd90f53f8db0629fc9b06ce;
mem[694] = 144'h0531f2ee003805ba084d011d07e0fde4fa39;
mem[695] = 144'hf93ef88a0549f22608c4fa090614fac7f27f;
mem[696] = 144'h00ea08c5fe2dfdbef9ddfd2e01bf05ac0d45;
mem[697] = 144'hfee40c41f205f7b900d9f5ec0a06f84bf974;
mem[698] = 144'hfc3ef3cf07f7f2cd0779027e0cf006d7f45e;
mem[699] = 144'hf0e8fcd40bf8f18704d604870c2ef0f8f9cc;
mem[700] = 144'h0595f1ec0c74058a0d5ffa9e02a00b0e0d89;
mem[701] = 144'hfc02f6d9fc2c0c350075f6da0894f4adf739;
mem[702] = 144'h06530ed2f967f4a10bd1f69bfacb0f52f1a2;
mem[703] = 144'h067509f2075df2e109a90845ff8d031df4bb;
mem[704] = 144'h0572fb9ff41e00ca05bf0baa00c607c0f73b;
mem[705] = 144'h073e0511ffca0a7afcbff848f0fa05e00dce;
mem[706] = 144'h00eff863fcf3fac40969f950f241030b0ced;
mem[707] = 144'hfb2d00ccf5c3f958fbb3079cfe820919f1c2;
mem[708] = 144'h08b20777f73b02f4093601a0f0210842ff7a;
mem[709] = 144'hfd81fb6e0a0e0702092ef158fe24f258f565;
mem[710] = 144'h03b6fa510bccf7eaf03c00260245094604ca;
mem[711] = 144'h0399f01df7d5fd5909270d9ff2c307e90ad1;
mem[712] = 144'hf5a6f630011a02c4f671018eff1f0dbf0f68;
mem[713] = 144'hfaf2f9590ea2f7dc0b03f6ed08340beefc03;
mem[714] = 144'h00ccefe1f89801f5052e005003b9f664fac0;
mem[715] = 144'hf2a4fc120ba20328f2330f00f138f6f0052d;
mem[716] = 144'hf8c80504f75af79cf4c1f627f928006605bf;
mem[717] = 144'h038e004dfd0a09a1fe7800370aeafdc70560;
mem[718] = 144'h0a59fe2b0bca0a4604d8006bf07e0a110ea1;
mem[719] = 144'h05930b9306ebf441f22ef766fa2806720f29;
mem[720] = 144'hefc80e1ef1150a1804ba0c270db90d4ff8be;
mem[721] = 144'hf3adf6dff7b50c8bf03a0f36fd330081f86d;
mem[722] = 144'h0c5006fe044cf8a00a09f684fe1a019e04b4;
mem[723] = 144'hf6ea0789ff21faf7f463f48d0861f8f3f5ad;
mem[724] = 144'h0f1c0f2b06590a64f63ef25a0f1205430088;
mem[725] = 144'h03660ded0e51f3ee0f5efaacf8350028f393;
mem[726] = 144'h0dfc0a5cff72f374f5aa0d9505b807c2f524;
mem[727] = 144'h01ea099bf6b706cc00c7009eff45f97c01b1;
mem[728] = 144'hf505f27c071ef360098c0f850ca60b040504;
mem[729] = 144'hf6faf811f570f45504d2fdc3fcb7f615f858;
mem[730] = 144'hf84e05cff041f16cf5bc0151fe530c550deb;
mem[731] = 144'h0f760a0c0d3cf699f63302ecf9470e2500f2;
mem[732] = 144'hf3e2fe94fbaf0601006c0f67070b0acaf7a3;
mem[733] = 144'h042a0c26048cf018f964f931058907bef9a0;
mem[734] = 144'hfae4f0ddf4cb0401072bf6cc034806adfb32;
mem[735] = 144'h0040f6cf0403f1370d51f6b7fe670b6e0cc2;
mem[736] = 144'h053106d7fbd609ca054d093ceff100b30e14;
mem[737] = 144'hf432f65df1870c99ff34073609c2068dff45;
mem[738] = 144'hfdf80b7403a1071ef679082a010d0b58f3ee;
mem[739] = 144'hf36cf3a2fd1a01e4fa64f7e1f7e0041d056d;
mem[740] = 144'h022ef96af1dc057404e7f591fc9f0bcafce2;
mem[741] = 144'hf427078909840c2c01ddf5900243ff2bf188;
mem[742] = 144'hff09fe850bfd0e8ef7f2ff3205680bc8fdfd;
mem[743] = 144'h08d8f6fc0c52f261fd200e1e05b50a0cf328;
mem[744] = 144'h0ea20bb2f58609430c7c0aa50f5a0a29f3ec;
mem[745] = 144'h065ef4e003190d3201090e95f47ff985f414;
mem[746] = 144'hfe3af3780af6f7e50ad8effa0193f4d701aa;
mem[747] = 144'h06920e7d0286fc0efdeaf8930d41f24509ef;
mem[748] = 144'h0f1e078d0c75ff78055f0bbff2ccf84ffa9c;
mem[749] = 144'h08bef7990fa909e202e007df040ff9ab0344;
mem[750] = 144'hfc0bf18a0abef1e3f8760880088af1bf0057;
mem[751] = 144'h0317ff9cf13403d8095701a1f48902cef7ef;
mem[752] = 144'h0eff0b34fe16022f0e420315f46efb9d0b57;
mem[753] = 144'h053700f2049f02080f57058f0c510511043a;
mem[754] = 144'hf7420b29f5e90820f9a5f8d8048ef710f46d;
mem[755] = 144'hf327fb9ffc2ff23cff730517fef0f75df971;
mem[756] = 144'h07500e42fe3bff470d5f0591f2b40cb60835;
mem[757] = 144'h092c03f7027c0dc6f687059a0627fa67fcc3;
mem[758] = 144'hfc0af37902e8f6830799f7090a68fe78f476;
mem[759] = 144'hf7370440091d02410d70f713fc7600730190;
mem[760] = 144'h0c370b6bf80ff6a9f9730051f380046d05ab;
mem[761] = 144'hf94402940342f35e0253ff110733fe0a0a41;
mem[762] = 144'hf72afa28fab30e03f66103a90e36078af095;
mem[763] = 144'h015cf782f9280ce4f6710d4807f30504033f;
mem[764] = 144'h0824fea8f7dbf61ffca60538f16508aaf591;
mem[765] = 144'h0152fb1af22af39e0035f1f7ffd3fad1f5fe;
mem[766] = 144'h00a1f8b20310fae5f36e0d0ef02e0b0afc02;
mem[767] = 144'hf77af1dcf391f8e0fb40f78906eefd230a1e;
mem[768] = 144'hff16fda5f8f1098cefee07fd0baa0e0300bd;
mem[769] = 144'h07560570f5e102ff016a0032fb10ff3701ec;
mem[770] = 144'hf4a6f655052cffacf3b0090d02f50170043c;
mem[771] = 144'hfbcbf3360c6ff6120a97f22e0bcaf92905d7;
mem[772] = 144'hf1b904d5eff2f87af284f93a07db0a1a0879;
mem[773] = 144'hf631087dfaa803c207360e0208d107600a79;
mem[774] = 144'h01d6f1af0cdc060affc7fadef7660cd30145;
mem[775] = 144'h08ddff7ef5fc0b7cf371fa260dbd09f2f9d1;
mem[776] = 144'hfb6cfb1d0a2e06d70dccf933f9140ef2051d;
mem[777] = 144'h033b0698f14807e5047a07f20be9f4560e7b;
mem[778] = 144'hfd5ff844fcc10b040048fd53eec4f26a02c1;
mem[779] = 144'h0426fdeb0873f6c30582ff3d0ba8efe4f4ea;
mem[780] = 144'h064109b6065b0052f70ef982f1a407d2f9fc;
mem[781] = 144'hf83ef6540682020cefe3fe5ef6e808e5fcff;
mem[782] = 144'hfd9b01930c4efebb0378f028f6eaf98df855;
mem[783] = 144'h046ef510f687fe0afd40fd56f4cf0261f0a1;
mem[784] = 144'hfbf2f4eeefe3f147f8abf7d0f6e1fcc90cca;
mem[785] = 144'h09a8026ef95804cbf8cb0cee0f60ffdef617;
mem[786] = 144'h02d50b3df9f7f813f3a90a960db2064efee5;
mem[787] = 144'h00c5fd04f600feba0ff80f71fafe05fdf445;
mem[788] = 144'hf1b6f120fa89f86c027005b6f335fe7df061;
mem[789] = 144'hf063f9b706c8ffecf38cf2c9fc0cfaf101bd;
mem[790] = 144'h0a2608bb0fe7f98f0e74f2ed00f3f43bfb67;
mem[791] = 144'hfa4bf0a1f73005890d43f531088e06f50eaa;
mem[792] = 144'h0943ff8b0187f768f112015c0eb8ffb10457;
mem[793] = 144'h0cf0f26d0535f7d80fb10d0cf1fa0d530860;
mem[794] = 144'h099307e9f50c039cf845fe6204d9092afe25;
mem[795] = 144'h0890fe1e0b6c09a703c3fe67f5abfd7cf1f9;
mem[796] = 144'hff06f8d6f505040cf69e00ab05ecf72ff908;
mem[797] = 144'hf2c406160c60f3100a72f7f3feacf65bfb6c;
mem[798] = 144'hf7c5097afac90964015efd3007e8070ef67c;
mem[799] = 144'h0de7f45bf6bef54ef160074ff0330b560be9;
mem[800] = 144'h020aff9f06f1f118017e0f5dfbe6f0a9047e;
mem[801] = 144'h00f6fec409e5fd84fd6ff18af0460377f6e1;
mem[802] = 144'hfcdd01e30e3d0af400b90f29f337f196f6ab;
mem[803] = 144'hf4fafa59fc720614f4ae09b90fcef88e0129;
mem[804] = 144'hf09ffed6fcf2055e0f38ff1dfbf5fbf9f53d;
mem[805] = 144'h04f70d7cfee7024bfb01ffd3f411f021fda1;
mem[806] = 144'h078903c0f9ca08280c370d46fd21fea80872;
mem[807] = 144'h0858fd75f89c0c71fa5100baf1a20fbd0d79;
mem[808] = 144'hfc96fc09fdb5fdd7088208bf0e4907a7f5f8;
mem[809] = 144'hf64c089d07ac096e011d0b18f7f902d9fd91;
mem[810] = 144'h024dfc51f731fe3c07930e1e057605ed0590;
mem[811] = 144'hefc6f4adef76ff6aef48ff7cfb0a068d0f1e;
mem[812] = 144'hf3d805e3f08afbfc0d7e0d05043203b509f5;
mem[813] = 144'hf4580b120d5befbe0236f60b0851fc75f4b9;
mem[814] = 144'hfef10f06f3f3fc950a25f652f35507410489;
mem[815] = 144'h0f56f3d20d9308040ebbf1a804530cceef6b;
mem[816] = 144'h0a55fe21f6a9fdd50b04087cf3c2ff3b05d5;
mem[817] = 144'h0366048a0c0b0b76f9f7f9bdf58c08d80382;
mem[818] = 144'hf3f4fd24f18bf8fc0dc309dcf9c9f7d9f0f0;
mem[819] = 144'h06160b18011b0c95fb4d039e070302adf922;
mem[820] = 144'hf3580ca703acfc36009afa1605fe089f0584;
mem[821] = 144'h06510b6cf5a8f9930c90f9e50197f547f82e;
mem[822] = 144'h07e10d7f0407f0f0fda90729fdef0492feeb;
mem[823] = 144'hffe00ac4031c04140bb50cb1f796f6650d98;
mem[824] = 144'h0760fbb308940ddb03fff17ff8e306dafe57;
mem[825] = 144'h080afa21f26b0aeef19fef5cfb370e9800b7;
mem[826] = 144'hf5ec06a607b50771f696f0db0a0bf8b3f56c;
mem[827] = 144'h0e2307f1fa3f0ab303a502d60074f9f20307;
mem[828] = 144'hfad904ca05610b3df6d9f7dc09200c8b0a60;
mem[829] = 144'h0db6ef95fb68fdd50d6af550fd58fa5d00b1;
mem[830] = 144'h005606d9042af3f80c8afe120a49019f04ad;
mem[831] = 144'hfc6cf656f7aaf984f8a10ce70c57ffdaf427;
mem[832] = 144'hf829fee9feeef280f3eff3ac0ca4f61c0bef;
mem[833] = 144'hfab0fbdfff320ebf034efe640d4bf6c7fc4f;
mem[834] = 144'hfc36f5eeff750ac7f5730c5afed90807f651;
mem[835] = 144'h0986fc37081af383093bf680f9690ea0fddc;
mem[836] = 144'h0f54ffaef732f5eefdae0bc500ecfd47fc0d;
mem[837] = 144'h016d09be01970009ff9ffa9e0f59f6e7f1dd;
mem[838] = 144'h035bfa240644f6650638f66b0313fca40deb;
mem[839] = 144'h02fa00030efcf8370d6703620ae104a2f13c;
mem[840] = 144'h089f0080f9ea0f5602d0fc7afa1903e7f569;
mem[841] = 144'h00e3078af15f08abf760ff0aef250f42f931;
mem[842] = 144'hff47f46f0b8cfa2bf7d20c280e3a0e260f85;
mem[843] = 144'h05b906c5f5ebf2e10a83f2a3f1fdf90af260;
mem[844] = 144'h0a6808befdb704e50053fdfaf79cf360f984;
mem[845] = 144'hf29c0a5f0d0607080f61f791fb33fbfffa03;
mem[846] = 144'hfd52013cf1a7005e00a80249f3cb061cfdbb;
mem[847] = 144'h06a603120b4404a105580784fddd0a620743;
mem[848] = 144'hffe1f66ff0e3fd09065e0654f3bbf9a2fd5d;
mem[849] = 144'h0603f1d804050acd06e3f1c0fb0109dd05da;
mem[850] = 144'hf0740a430f89f5c90b1600980a4cf9790a78;
mem[851] = 144'h069bf504f55a079ef9bffca00a72f8eaf71a;
mem[852] = 144'h0c5c004e07600deff54a0cc80fa2fc020ade;
mem[853] = 144'hef180c4bfe2af102fd7b04d3099c04d00e2f;
mem[854] = 144'h097207dcf4e4066afa6c0333018009fe07c6;
mem[855] = 144'h04adfaec06abf20bf2cc0307f87206ee0f45;
mem[856] = 144'hffef0dccf9ebf29106a60500fb5bf6340b83;
mem[857] = 144'hfe68099707b70ca5f7b6f56a03a10b520293;
mem[858] = 144'h0b75fb0cf27ff7440e5df58104ecfab5f298;
mem[859] = 144'hf406fe190aaef2ff0da70737fc82fd74fbe3;
mem[860] = 144'hfe38fe28057dfee70156f2e5f4dd0ae70479;
mem[861] = 144'h017df6d2f249037b0c21faf3f225f94d0375;
mem[862] = 144'hf71ff69f0eea0107090e085003270ba5f3dc;
mem[863] = 144'hf0610f62fdc0fb48f4c7f8e5f6acefa9f5bd;
mem[864] = 144'h019afa3d06a7fd6a090600ce05fa002d00f2;
mem[865] = 144'hf04a00b20d6c05d1f64808aa00b8fa6908e7;
mem[866] = 144'hf4d5f737fae604effbc5f7c9fa62f70e0e1a;
mem[867] = 144'h01c9f3bd0581011807f1fd8706baf01d0127;
mem[868] = 144'h0ad8fb81fb82055f0399f74e015af9f0f5e1;
mem[869] = 144'h0cf8f9ab082903550560038209f9f1b1054e;
mem[870] = 144'h0826f0e9f8a507eefdcdfce4ffc7fe53047a;
mem[871] = 144'hf4a0f104fa5ff7630943fed3efeaf8d806e0;
mem[872] = 144'h0226f39a099307bff90bffbb05340279fc23;
mem[873] = 144'hf7a2f4d9fc0bf6d5fe4c0683fd43f6a5fec4;
mem[874] = 144'h084d0a02f9e6f10f0376ff6f0cf3fb970c1f;
mem[875] = 144'h07e9fe1800b1fe5d0705f335f4ebfadff346;
mem[876] = 144'h01f3090b0e46f5f1f45b01bdfbdbf59c0ae2;
mem[877] = 144'hf964efecf83ef28ff0e90156fa1c0d6501d9;
mem[878] = 144'hf680fccffdd7f4aafafb0cec0e79076606ac;
mem[879] = 144'h0f2100cf0080f47cfa63f650f082fd47f390;
mem[880] = 144'h0ee20b56ff8d05bcf0cafbeaf7fe0e74ffa6;
mem[881] = 144'hf9350bab0efffc6bfa670593f5fefd4409ee;
mem[882] = 144'hf4a10e73f152f082f15afcc6fd19f0790ca3;
mem[883] = 144'hfec70cb4055ef03bf314ffca0932fb5effba;
mem[884] = 144'h0e22079fefea0d82fb82fbe0ffc20ba0f0ed;
mem[885] = 144'hfe0c045e011af185f5c2043ef0930d27fc9b;
mem[886] = 144'h0d8dfcdb0611f399efccf9c8064dfd7506aa;
mem[887] = 144'h0997f1c1f3020588f2d5016303a60364ff1e;
mem[888] = 144'h02300519f7e0f37fefa9f71ffc60023e0c8f;
mem[889] = 144'h0356fc10fc5a020b0301032a0c14f0bf074d;
mem[890] = 144'hfe6106f4f69308cbf43b0ce505b408d70d0e;
mem[891] = 144'h02f309080ba2fd680c60f9fdfc0706c0fece;
mem[892] = 144'hf533fcf60b3dfca5fa1402ff0eb8f7650baf;
mem[893] = 144'h0d2dffe0086806d8f9e2f9ebf4e40318f2de;
mem[894] = 144'h02e70ec8f89efbfe0f77009902b7f6da0bdb;
mem[895] = 144'hf443efc4fa3afde9f8e5f881f71e0680f3e6;
mem[896] = 144'h0457fb980e3ef2b80eaf00620578f681fdac;
mem[897] = 144'h089df887064cfc53fe01f3bbf41df1830634;
mem[898] = 144'hf1c10f5ffff5f425fe3c0c17f1dcf5cd05a7;
mem[899] = 144'hf4b80d8702c70040041af8e70633f0de082f;
mem[900] = 144'hf55bf052f829f1ed0f5e068df72bf2ccfc97;
mem[901] = 144'hf8eff94104f402060446073ffcc701fbfd07;
mem[902] = 144'hf71c0bf3055e019a00e907c40b29f2adf08e;
mem[903] = 144'hf85c04a7ffc907030f54072d0543f31afcf5;
mem[904] = 144'h04d2effe04410eadf87df7e00c28f5c30ccc;
mem[905] = 144'h0aeff77d084ff6f402defb520694f8f30a5d;
mem[906] = 144'h003c0a93f6f90ec8f13d003f0e3a051d0bca;
mem[907] = 144'h0aa0030507b4071207260375f79a0373f196;
mem[908] = 144'h0cbb00b70d60f86c0032f4d4f9070f97f946;
mem[909] = 144'hf8e1fd17f46df44801f30fb30f4d06230285;
mem[910] = 144'h0d3af536f25efacbf50b0e9df8a40eabf0fd;
mem[911] = 144'h0db30164f376091afa340346f5cb0d7001db;
mem[912] = 144'hf196f407fbc702570200083af93706570064;
mem[913] = 144'h0627f8b2ff070a19ff8300f40106f4b8f5b7;
mem[914] = 144'hfa060ba40c60038c0778fc810d09fc92f57f;
mem[915] = 144'hfc510745f0960d7efb6007f00fd5080e02e7;
mem[916] = 144'h0aa5fb05f11b01970a82fb4b0a6ff60ff5b8;
mem[917] = 144'hf6870337027ffff9fcfdfe1a01b7f7d5f6f2;
mem[918] = 144'hfdbf0f260a18056afe80f6b60f7203620af0;
mem[919] = 144'hf5db090ffb9e0ce0f40b0870f257fb36ff2f;
mem[920] = 144'hf9faf270fa6bf36f0601fca50620fc4df4d9;
mem[921] = 144'h0997fc3df39e092ef9afff1906f10afb02cc;
mem[922] = 144'h066af03cfe640be007fc0c04f89d0491f09a;
mem[923] = 144'h08b10810050c07e109d4f7d90dab087efe67;
mem[924] = 144'hf6410d100e28f5a2058c08130aa20d1401c6;
mem[925] = 144'h00390a1ffe09f615fcc704b20d97fbfcfc3a;
mem[926] = 144'hfb60038d0a96f8d20120078000390c35f97d;
mem[927] = 144'h078d0d19079ffac8f3ccffec0ecf0e33fb21;
mem[928] = 144'h019607c3fed800b6fae206d6021a0b390d79;
mem[929] = 144'h06d80ee0063af38102530d5a0b6e09fb0a13;
mem[930] = 144'h08c1fec8019803db07890bd609d9f469fe3b;
mem[931] = 144'h03cdfd37f609f2eb02dc0b22fbd2010b042b;
mem[932] = 144'hf628f032f8c206110c93f515f109f5fa06c0;
mem[933] = 144'hf7c001f5fea7f22100c8017003010153005d;
mem[934] = 144'hfc8cf4c70c0f0a5dfa580758f80def660570;
mem[935] = 144'h0b8a0dc3f2710541f538fe27fb91f5980438;
mem[936] = 144'hfed40623f8daf5bcef0cff83f1a1089d0560;
mem[937] = 144'h093efcd2f65a0416f6bd04e4f168f975f76b;
mem[938] = 144'h0e29fecff167eee1f1770ce1096c08700cea;
mem[939] = 144'hfdf30833f9100793fe1d03270d8aefddfe8c;
mem[940] = 144'h0a7e0a79f95bf5cff5bdef43ef81f1befefc;
mem[941] = 144'hf401016efc89f8cbf9960213fb82f3cbfd89;
mem[942] = 144'hf2bf0284084c0428004e0aa6f2fe067e0df6;
mem[943] = 144'h0d0f0b3c0d390c2906deef35ef910897f2ca;
mem[944] = 144'h0188f5c9fae1ff0f0c5ef3e9f716057bf6ba;
mem[945] = 144'h0c7a087201d400f9fe04fe27f77b025bf821;
mem[946] = 144'hf0caefeb0de7f2880c5ffc7ef1d30623fb55;
mem[947] = 144'h0802040a02f2028b0c06041104370f390db7;
mem[948] = 144'h0cfdf431f79f000504a8ff21fba0f3fbfa69;
mem[949] = 144'h08940e580a97081ef6cc098bf746fce4f612;
mem[950] = 144'hf444036aff5d07c60da90327f992f74efa3e;
mem[951] = 144'hff93f17ffa9dff6306380d1aef180c470ff9;
mem[952] = 144'hfa2cf8c304600984fb89f64cf0b7fe380699;
mem[953] = 144'h0556fd0ff2c6061804c9f695f0490cc5fa12;
mem[954] = 144'hf53e016a06600e83f4b9f37b070afcf10b41;
mem[955] = 144'h0b970c8afb160a5b0bf1f8eb0abff1dc09d5;
mem[956] = 144'hfc2cf530f8120d5bf8f5fe48efbf05b50e4e;
mem[957] = 144'h0e3efe390e92fbceffa004cd09c50c3501b5;
mem[958] = 144'h04f3f4960bb3f92f0dd6f3ddef6807c80756;
mem[959] = 144'h029502e606c6fed3030cfaa40cf80733fdaf;
mem[960] = 144'hfe8705440b830bf7fe24020f08af0a16f2aa;
mem[961] = 144'hf34ef9190c920f76f50509c60776f3def594;
mem[962] = 144'hf705ffdd045e0590f9a3fdff09fd02c10f26;
mem[963] = 144'h0388f4c101770e3709d80f0d03eb03ca0262;
mem[964] = 144'hfed90b5dfb55fb630c66f11d011409f8f1a2;
mem[965] = 144'h00a90e7e055306eeffaaf345fcc4f0ba04e4;
mem[966] = 144'h0584037ffe0bf0e2f532fcce0b6d08850610;
mem[967] = 144'h03aff833fa13f1820280027a0568f89c0ae8;
mem[968] = 144'hfae90f1400fa04a10a2befa2fae70897f5c6;
mem[969] = 144'hf10cf7430c97000f00b4fb65f7bbf4a0f517;
mem[970] = 144'hf9bf0220007c0db1fefcf623ffc6f05e09e7;
mem[971] = 144'hf4f2fb8cf4e906eb0138fc0cefdbf988fd8d;
mem[972] = 144'hf6dafd260ea7f70af824f5a7066206ba056d;
mem[973] = 144'h0f63069cf844fb32fd81feacf6ad061b0c60;
mem[974] = 144'h05ef0549f03002880adc08e4056903420442;
mem[975] = 144'hfe820ce3fff9073d0a7ff90a02520498fcec;
mem[976] = 144'h091f0acbf7b5fdef003ef4ff04d3f470fd86;
mem[977] = 144'h03baf98af34e0a4205b3f7bd0ea40704f819;
mem[978] = 144'h0256f1e1084bf5b7f9def95df887f7dafd5a;
mem[979] = 144'h08570592fdfc0df407cff0fff0300a2f0e70;
mem[980] = 144'h0811f302fb1b000dfe9b05a4032af662f2dc;
mem[981] = 144'h0bf9fb280d31fa8506030beafdcdf302f059;
mem[982] = 144'h02cc0af1f5b1f25ffc44fe25fbdff4fe0b30;
mem[983] = 144'h0f13f1b60c7a05690845f7c20326fe7b06a9;
mem[984] = 144'hf4eff3840abd090ef6e8f105f9d7f6baf0be;
mem[985] = 144'hfbeefad30c4b0116f69cfbf1f68002fd0b31;
mem[986] = 144'hf00f018b088dfe64f2c1070f043cf7f60326;
mem[987] = 144'h06650e0d080efae40edff2fa0e93faedfc6e;
mem[988] = 144'hf643fe5902f6fc66f48ffb4c0c6309c80624;
mem[989] = 144'h00f8073503c806a3f8910eb4fd25fdacfdc9;
mem[990] = 144'hf02a011909ac08ab0402f17b07acf6a1f06b;
mem[991] = 144'h01daf236fa59fb1a07bc0e830495fb2c0118;
mem[992] = 144'hf74d08f4f5030c72f2e7feacf9a30540f1d5;
mem[993] = 144'h04bf0fda022f0a85f8f203df006803b506d6;
mem[994] = 144'h0ae2fd1d0d3ef01100f901f0055b0a440d4c;
mem[995] = 144'hfec3f8dbfd250505fffc0014f6c2f30ef4a2;
mem[996] = 144'hfb610ac9f74bf995f9e30c3bf684f984f8dd;
mem[997] = 144'h07e4f4b0f7150cdf0bc6f10e0c9b0b3bf704;
mem[998] = 144'hefff08f30bf10a720e5f0092f5e8f30ffd68;
mem[999] = 144'hfa380302fd8cf84efb7e063d01790b13f80a;
mem[1000] = 144'hf65cf0e9f3aff98f051606990acb07e40906;
mem[1001] = 144'h00ddf1f9f54f07b4fa3defbbf41af994ffa6;
mem[1002] = 144'hfcddf1880557fa15f21e0720fce7f6b60ea5;
mem[1003] = 144'h00aef282f25b0b39f1e4f45cf01806d2ffcf;
mem[1004] = 144'hf33503aef4ba0288f1e6ef39f0f8fd0c0ee8;
mem[1005] = 144'hfdf7f9d40c370b3301f70e8e0d4b01e2042f;
mem[1006] = 144'hfb9df4e30bcefb970d5a0aac0b040c3b0725;
mem[1007] = 144'hfc5c008404e7f26c097cfe35fe05f3a7fc4e;
mem[1008] = 144'h0305f3040e970050f725f0800624ffcf0ca6;
mem[1009] = 144'h0132f9940da4fe5c059c017cf784063df3c9;
mem[1010] = 144'hfbc3ff8a01810f15f711fad60cb20553f4c6;
mem[1011] = 144'hf5c1f0370ef3f2fbfa40f827fab9f55cf1e2;
mem[1012] = 144'h0caaf1ce0915f15502510556f3bffd5eff32;
mem[1013] = 144'hfa74ffa3fb8cff65ff790e43f4f8fe31f9c6;
mem[1014] = 144'hfd1fff900b7f05b2fb88078d0508038b006c;
mem[1015] = 144'h06adfeb60636f9e6f31603b8f4c0f0c109a0;
mem[1016] = 144'hf175f9a2fdd301dc0c8a06ae0c44fd69089c;
mem[1017] = 144'hf7b1080b0e9bf4ca00c6f962ef39fd8e06d5;
mem[1018] = 144'hfaf50bcf03f1fd8706e30346ef520eaeff12;
mem[1019] = 144'h042ff8f9fe83fce30b03fca30c0d05ca0c04;
mem[1020] = 144'hf4a4f9c2fbd70380fa200b71f45102d9f9a9;
mem[1021] = 144'h0dcd0969f6e4fefa0c68f5b1f0cb0f8d0bb3;
mem[1022] = 144'h07a805c503e40b75f376051ff5740ea9057c;
mem[1023] = 144'h09f6f66a07c0f9fef7690102081ef940f215;
mem[1024] = 144'hf716fe11f761fe21fc8806d70560f772f1d6;
mem[1025] = 144'h0e970872fe27f969fb750d960c5cfe990b57;
mem[1026] = 144'hf5d1fbcefeb8f5f5fea600d5ff8c09ecf8c4;
mem[1027] = 144'h00cd0ad2f3e406c0f2b5f2ae0e6cf86cf600;
mem[1028] = 144'hf73b0724f7f20427fd1c0ec4faa707490413;
mem[1029] = 144'hfc8809e90724f40d014a01ae03ce0ed8f177;
mem[1030] = 144'hffb1040302d8f05a08880041fb96f8c7f4ce;
mem[1031] = 144'hf97103b1fa65f2b402b905cdff1cfd09f189;
mem[1032] = 144'hf6aef1760cd1f744002d0b9bf06af00ef319;
mem[1033] = 144'h0812fc20fdb80105f3a4efdf0689f5fdffcf;
mem[1034] = 144'hf833f5630e3d0776fb78f6ee0ea701310791;
mem[1035] = 144'h0a89093af84ffe0ffc2fffe304e5fef607ff;
mem[1036] = 144'h08180aa5fc150033090801280ae7fbc4f7ca;
mem[1037] = 144'hfb860d00f7d10037f007facc03b201bbfa63;
mem[1038] = 144'h0007fe66f542fd7b09bafe93fdeefee5f463;
mem[1039] = 144'hf3ff0f43fdf4023807ef06a504e40b31efc1;
mem[1040] = 144'h01d2efdd06a3fd71f97700b9f1c7fa1c05e9;
mem[1041] = 144'h0397f038fb95f96b0e93f161f8800bf70308;
mem[1042] = 144'h08e309c40466fa38070805250844022e0e48;
mem[1043] = 144'h0fbb0eeefccc0b680736f727028df7ebfd9d;
mem[1044] = 144'h0bfdf551f8a30d09ffd2fa4303020c10f5e0;
mem[1045] = 144'hf23e0e62fba6f666f6d80a18fa3d0e54efeb;
mem[1046] = 144'h01d0097f0cf4f8c1f5910e33f991f6aef788;
mem[1047] = 144'hf13ff953fa980a11f8daf750f252f961f799;
mem[1048] = 144'hf5e2f5350107fcb20293f14bf6860218f1f1;
mem[1049] = 144'h02fbf921fcc9fa84059cfd10f08af34efd82;
mem[1050] = 144'h009c03f8039d0919f6650009ff4b0d080c15;
mem[1051] = 144'h00e90b3b0caaf7be0bd1fa7ff5430b35ff4b;
mem[1052] = 144'h060807690b2d0c82f811f1050e7dfe8e0665;
mem[1053] = 144'hf2170e7ff991f96df9e20be0ffc9fe9d0041;
mem[1054] = 144'h045dfae5f2d20299fc3507f4f8da0b800af1;
mem[1055] = 144'h0edb096d00cef3f7f2ba082f08fef362f12a;
mem[1056] = 144'hf4f502e00eec006d0de1094bf7b60128f3bc;
mem[1057] = 144'h0f26062efd1dfe54f1dff96af0a1fed5fa4d;
mem[1058] = 144'hf605f6fefebf0e280dba0fbf041f0dbffe0d;
mem[1059] = 144'hf29b06ac05bdf22e0b7008ab0f4df96cfe6c;
mem[1060] = 144'h021af555effc06e808f50cdb03a40f1df289;
mem[1061] = 144'hf5c8067ff159ffa50eac0858f9470558f24e;
mem[1062] = 144'hf5fd0158048607d2fa7cf985023cf94f0cf1;
mem[1063] = 144'hf6a502420c7bf903fb3900defb86fdcdf446;
mem[1064] = 144'hf57a09730aa108bf06cbf08b040ff8a6f372;
mem[1065] = 144'hef89030af9b9046d0731f2f4fcb40985f74e;
mem[1066] = 144'hf4c1fdd403760f1b0d7ef0a1f856025df1cf;
mem[1067] = 144'hf2effa5aefc604d708ac00ac03b00331f178;
mem[1068] = 144'h0f97f0b101edf7f1055401c0fb990a55f440;
mem[1069] = 144'hf7440287f4040270006401a7f565fa50f3fe;
mem[1070] = 144'h00aefeba0b9005a40ce5fec40e770d460193;
mem[1071] = 144'h006201f7f768f82c0cdf002cfbbefd1cf968;
mem[1072] = 144'hf20201a8f5acf6b1f172f3a406d70394f227;
mem[1073] = 144'hf215f8def69af01df0a7f06c09a30240002c;
mem[1074] = 144'h01250265000004700ef605a500a20cd4035e;
mem[1075] = 144'h0bcef316023e03e800fcf385f6f304440653;
mem[1076] = 144'hf4ca0c080901f53602fa0edd008302fd0070;
mem[1077] = 144'h03eef2b50d200f730cfa03ecf437fda9f66a;
mem[1078] = 144'h05def506f923f744072efa910b11fc5b0990;
mem[1079] = 144'h03cf099ff8370c060f600996f9ca0ced01a2;
mem[1080] = 144'h0b12f57108c604600086fd3ef771f1eef7ae;
mem[1081] = 144'h0690f0edff620bee0940fc4407350aa2082c;
mem[1082] = 144'h01b4fc3b019c0cdff9ccfdbb0cd00afd0406;
mem[1083] = 144'hf30ff531ff27fce70a5c01d60e2e07d7f5b7;
mem[1084] = 144'h0eb9f7d309780b7dfc13fd39f51807e20092;
mem[1085] = 144'h0b670e0ff2fdf8880f0f0e560aa4f9880491;
mem[1086] = 144'h070e06d1f2c3025f038cf88c085df228f7e2;
mem[1087] = 144'hf34df8fbf6bcff87fb1d0a97f2120afbf8e6;
mem[1088] = 144'h04abfb60f71b0cc3fa08f337fb5901b10b91;
mem[1089] = 144'hf63e0523f247f61af300f228f9b202b20f77;
mem[1090] = {16'hf3b3, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1091] = {16'hf0bd, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1092] = {16'h0d7e, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1093] = {16'h0860, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1094] = {16'hf166, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1095] = {16'h038f, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1096] = {16'h01b4, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1097] = {16'h0010, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1098] = {16'h089e, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1099] = {16'h0399, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule