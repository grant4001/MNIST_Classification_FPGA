`timescale 1ns/1ns

module wt_mem2 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h110be0b80aee1b0814720fd10682191c0e53;
mem[1] = 144'he48a113f03bbe33b1b69fde001aee813e0c1;
mem[2] = 144'hef65e86904edf9d81c61e422e62e1d20eefc;
mem[3] = 144'hee31f467e579e784fb26f0ccf2fd00811344;
mem[4] = 144'h1309e87b1da413720967081f0d71006311bd;
mem[5] = 144'hf89ef29714c30550077f1ee5f01ef0fb0ebf;
mem[6] = 144'h188afa59f49adebdfd021253fc361010fda8;
mem[7] = 144'hf7691168ec4a10dd1bb4e8e3082f1e410c90;
mem[8] = 144'h0b12ff2915b5ff47e94603d7eba5e36a1b45;
mem[9] = 144'h0426ed2ee6c308f91ca9e917fab0e541eaa7;
mem[10] = 144'he895e493fc44ed9bef85e0e81947e3771a06;
mem[11] = 144'h0f5d1e1ef774ef07177cf7a10f0ae5850bd8;
mem[12] = 144'heac5f430185cec8fedfb0c93f452f0660394;
mem[13] = 144'h0cf9029e13cae9d40b810fe91d05e257e7b1;
mem[14] = 144'h0da3f86319a8f57d086013480916e0f00f21;
mem[15] = 144'hf3c40c641b030e77e09d1155121a15f7e2bb;
mem[16] = 144'h0082f54d1c600ced141be09e1dc30d98f668;
mem[17] = 144'hec83182e1b0e0e17054713390e32e487f24d;
mem[18] = 144'h163404edfe651889e9b4f00802bd19fe1abe;
mem[19] = 144'he48cfbe6074018cf14e61464e423f94018b8;
mem[20] = 144'he6e103e7172f0058e00e1b27e79710421ecd;
mem[21] = 144'he460e1ac1d8afbed1d1910cbeb20fb8fe078;
mem[22] = 144'h0c8b018319cbef8ff06df7e6df821abfdf79;
mem[23] = 144'he5c2e3e001e1f4940e74152000bc039f16f7;
mem[24] = 144'h1109fd05e4b1f85110f006c60c35f5a21c17;
mem[25] = 144'hf5650cee1d0f062ff82602bc19ba0f090290;
mem[26] = 144'h13831b7208e5e2a1f19b182e0d58e8df05a1;
mem[27] = 144'h105201d506871eb8e34916dcef0910701f40;
mem[28] = 144'h1139f349f29cf3c70459f8b8ecb9131b1586;
mem[29] = 144'h18cf1f8019b0ecb8f9c01fb4f94e0a2a09cd;
mem[30] = 144'hfc36f7b4151febbb1c8407ca118be1bc022d;
mem[31] = 144'he95414a1ff8705720e4409e9e4b21b4118f7;
mem[32] = 144'h1b701e831f741129f39ff420fb8f042df238;
mem[33] = 144'he5550f53144800b60194ec20f77a137de7ea;
mem[34] = 144'hedaa0f8a0bad014fe4e1e91afb3d16111727;
mem[35] = 144'h182b0fc2fddcfe06fdf2ffe1fbff1718ff32;
mem[36] = 144'h09700f95f0d3fcf90297194c1afff0aefca3;
mem[37] = 144'h162c14e41b3bfa201f710f4dfd9201890451;
mem[38] = 144'h0abae21f122f0e15f3b6fd801975dfc9f640;
mem[39] = 144'h1ffd02dc17e817501fd9e47ce25c00b21f2f;
mem[40] = 144'h1671f6edefe2f1241dd812af0a43e557e607;
mem[41] = 144'hf427129be35c0e84ed17134701030b670b6e;
mem[42] = 144'h0b3afcd7e261f7b5e2a11c6ae4df0ea50e81;
mem[43] = 144'h18adf2700ea9e15cf006ecf81605ff42edd8;
mem[44] = 144'h085619f11cfeeb82058e17d504b1147bed33;
mem[45] = 144'he36dea94f51bf7fc1a5ced121199f46d111a;
mem[46] = 144'hed3c12020896f81e1ced17edf0b4075d08df;
mem[47] = 144'hfc87170401ff008f0b5e1d2d01f21390e444;
mem[48] = 144'h0b160dcaeebce245fd2d093a00f704b7f7b6;
mem[49] = 144'hf247004af88912ff07160ea7e9230d0b18c9;
mem[50] = 144'h17b106e80a94ef41e97703201d4b140df0bb;
mem[51] = 144'h0b38f752ff880677eaf9f6b2f62a12e7119a;
mem[52] = 144'hf8940561f5c4e6a41d36efb4fb26ed32f25d;
mem[53] = 144'h011b17e3e16719cce54b13bbedf7fdc9eb78;
mem[54] = 144'he64ee3001606eb50e4771f0f0fc3ff29df5d;
mem[55] = 144'he711e8e0e0d1edde1871f82313e81b1ceabd;
mem[56] = 144'h089c0417f1ca05f8fb1b02dbffe4e4bd07fd;
mem[57] = 144'h1540f939f5de103ff6fe031d07cde5affd76;
mem[58] = 144'h189408c4e761e3030f8cf640e5951d7409b7;
mem[59] = 144'hfcb114bc1e20ef9f168a15d7136afde7e507;
mem[60] = 144'h0e540239fdad0b2d16ecfa2cf3dce30d19cf;
mem[61] = 144'he7dff12a0b6c051d0335e390f505eb8ce22d;
mem[62] = 144'hf6b51497f01be1b8f0980ac60059e35df624;
mem[63] = 144'h1461f52df5f70617fa59fd9b025512d1f78a;
mem[64] = 144'hf2b11ed70eddf818fcb7029ce776e64cf74f;
mem[65] = 144'he2171e74f887fb81016f189be2631a38f053;
mem[66] = 144'heba9ebe5014ff8ab0bd21910f762048b1ba2;
mem[67] = 144'h055df9a4f06512b40a0de231eab0e9d80657;
mem[68] = 144'h02dafb59f07cebcc1ba31a48191fe961f1e2;
mem[69] = 144'h1ad401310b2be4b10e06fc470d06ffcc1fa7;
mem[70] = 144'h040efe15fb69fd47e4e5146cf318e6eaeed7;
mem[71] = 144'h140d1c021f6f0799e10b08b4e354f3de05ef;
mem[72] = 144'h0138f1a513e1e578e3e1e8e81b99e611e7da;
mem[73] = 144'hf3adfb2203f80f3613580527f4ef134fe59d;
mem[74] = 144'he96d0f93ec4a02de03f217051ed7fcde1e7e;
mem[75] = 144'h02c60217eae61c980730efab0598faf7fa25;
mem[76] = 144'hf85deb431a670970fcecea36e7b50e31fa9f;
mem[77] = 144'h1e4c0506081ce25e088bfd09003605c10f69;
mem[78] = 144'h13a0e8040909e332edac169aeba9e7d6f39e;
mem[79] = 144'h06ad0727e407ff1c1d35ef20e8eb0ad3038f;
mem[80] = 144'hfedb00a6f9621f04f386fbd6e34aee330d03;
mem[81] = 144'h1bcef085e90a0076e2a00cb5e1def97804a6;
mem[82] = 144'he430f2a7ee6f17e7037e05830572fb03f995;
mem[83] = 144'hf3fdf7deea6b0191049b1b51fb371d8e1cba;
mem[84] = 144'h1033f1b71ce2ece505cf1cd705bcfe221a5d;
mem[85] = 144'hfee30cdb0e6b036119bb16ccee6216f1eb98;
mem[86] = 144'h12c3081cf366f2e0f688faaf0c09fd16e107;
mem[87] = 144'h1d5a1c1ffbf2e664f3d11a4f1e29073ceb16;
mem[88] = 144'h0d1901581dcf1f8c184a012d18b3115b17bf;
mem[89] = 144'hf4d11f2df68af94ee7d300a3e2521f0cfae8;
mem[90] = 144'hf485fb52ecd2ee26e7be190b05a0eeb7f6d7;
mem[91] = 144'he4e6e0ac06d7e4dbf42ee5e9f933efee1b14;
mem[92] = 144'h1b1f1777f9a2e273f19efbe4163f1037f025;
mem[93] = 144'he60e14d1f35e02121a8c1e180859102b03f2;
mem[94] = 144'hebabe146051bfdf5e12a0ead0c5614bd0018;
mem[95] = 144'he40f0f6be807041411911cf5eb970b8a08ba;
mem[96] = 144'h198d04e611a80706f2280867e1581537f8a5;
mem[97] = 144'h0826f115ee1d1b30078c12170c5a0db9f247;
mem[98] = 144'h0710fd8c044df339e0631c13ebbc0e27f848;
mem[99] = 144'h0b04fc5e080d063ff9bde2c8f4ec1815f9e0;
mem[100] = 144'h18251e98e2f5e8720068010b142c0ea1e3d3;
mem[101] = 144'he4b61235ee33facaec73ef6b1fb80619fdb4;
mem[102] = 144'he15bed7706371600f66b0e6107d9ed14fdfc;
mem[103] = 144'h108ffab6ea00f9c91ddc0767e0b10cf9ed68;
mem[104] = 144'he2ce136e1502fc1aff8afef10d5afb9e12d8;
mem[105] = 144'h1c71fbfce35cedea0ff808c100da0d4de3a4;
mem[106] = 144'hfeedf292fee21c80f0811049f4d8fe7317c1;
mem[107] = 144'h1c9319b01b5a04b206711aecf5571910eff9;
mem[108] = 144'h05840b9c0927e7e5efd2ec8de4140aa4ff7e;
mem[109] = 144'hee10f55effb3fee8e08114ee1ec10142e798;
mem[110] = 144'hfe35ecaa1196f096f2e4f52bf3201edb0d83;
mem[111] = 144'h061005281faef1af0dd81329e3fbe5b2fa09;
mem[112] = 144'h0d011123e09a0eb8135314bf0b2010c917c2;
mem[113] = 144'h03951683fc01e08e0b121322f02e055e14a9;
mem[114] = 144'h0ce6f6351fe2f99af270078fe4ece4ae05f1;
mem[115] = 144'hf969f857f01dedff1bccfe800453ff45e2a1;
mem[116] = 144'h19341dc1e157149fedfb0d410387f90d076c;
mem[117] = 144'hf5f1f0a8f906ee3f19991652e67d08f103c9;
mem[118] = 144'h0f28f994f16ef53ee8011600e6a0f25c0c90;
mem[119] = 144'hff82f32518d51e5a16781c6500bff2a41935;
mem[120] = 144'heeb31fe718c9f072f63bfd84fc49f8dd16cb;
mem[121] = 144'h17aa12bae142ea46ff081474138bf7db1fe3;
mem[122] = 144'h127af12bef53fdc216b413301f9df15ee53a;
mem[123] = 144'he0b4e4911370fe1401bee7a50b5dedb3e30e;
mem[124] = 144'hf6731347145ff2d0168f1710171c052e192c;
mem[125] = 144'he5a1e18a0f97ff0ae8b9ecdf11cd03ae0a36;
mem[126] = 144'h00f4f360ea741dd31084e561fc650dc51414;
mem[127] = 144'hf96901431072177e19e8f9c20544077e1e36;
mem[128] = 144'he7981c40fd8913a618f6ecd7f461e029e1d4;
mem[129] = 144'h0cb6e1c4ec53e297eac3ea55e2c01bdce1df;
mem[130] = 144'he725f45de8710123f81bf00ce9d60613e463;
mem[131] = 144'hee0de4abf0d9f759f738f8b714edfa10f2d3;
mem[132] = 144'h16c70e99e5a30f101cee131f1422e9fd0418;
mem[133] = 144'h029b1aa3f664fec914f0f7e5145ee3cd0a75;
mem[134] = 144'hf9bdebb20f801fbc002a0ab9f25bf6a90e20;
mem[135] = 144'h05f4e053ea88098be64df068e969ec271882;
mem[136] = 144'h153b0b9204f50ee314bd0fa3145b1b071535;
mem[137] = 144'h088b03121bbe068d2012129f1bf60d3cec70;
mem[138] = 144'h1d661f7feae8fdf3eb6ee88dfaf8f6a7183d;
mem[139] = 144'h08cff3bef495e3f8fca0ead10b7207ec1e8e;
mem[140] = 144'hf30b11a7016e0b9a05cdf1c9e3b40f690995;
mem[141] = 144'he5250b4e1026e1270e2bf81ae500f2b50b8b;
mem[142] = 144'h1b820e07f1f5108af8a40fb2f9ac0dfc1271;
mem[143] = 144'h1e1b0539e114068c04dcec17e46de984fdf3;
mem[144] = 144'hf3c6f40602b2e30a0a89fa5d0ceb1c36e126;
mem[145] = 144'hf0130208fe3312e40712143cf2f90b93fb78;
mem[146] = 144'he622fd6f1d19e3f5e960e69014ec172bed23;
mem[147] = 144'hef6afc2e1603f3061ca7022ef911e81ae20b;
mem[148] = 144'h0bba0e630124192ff72fecc8e274e9100ac5;
mem[149] = 144'h06baf4f715e1fff50a9fe1380be5ff0c13fb;
mem[150] = 144'h0d72051fee46f9c5fbba03a1067d0710fd6f;
mem[151] = 144'hf7dcf674e01d121be2a8ecaf026601d3ebe0;
mem[152] = 144'hfe46ec9f1ad6f8b71c97ffe716bd01f61ef7;
mem[153] = 144'h039e1706fc51e8cffde4fab9ff061382f137;
mem[154] = 144'hfe8cf4281bc2e4de1c8df193f0cef7461065;
mem[155] = 144'h1bd31a01f07ce6f9e7ae164ff7c0f777183f;
mem[156] = 144'hf5c2fb67e0a8093c036f0c6a1ee210431d72;
mem[157] = 144'h040aef53f3fde47c1381fba00dbf11f8eeb1;
mem[158] = 144'h036d015ee449e441f7cf0d9318efef0ceb2d;
mem[159] = 144'h0386026e187c0860fa8d0e48f8d51a9eeed0;
mem[160] = 144'h0bdd04ca05b009eb06ec1d73e030e956f51a;
mem[161] = 144'hf6e4ec5c005a0531149c0f51e5f61b7818f5;
mem[162] = 144'h0643ef19e7eeeecfe4c502f8f343fcb90e50;
mem[163] = 144'hf8ba06d1f96f1681e1ed1fe107c41b3a1753;
mem[164] = 144'hfa160947183cea38fd59e6d6164e19e4f578;
mem[165] = 144'h11b7eb4d1e5806960a070fb3f94ae84011b0;
mem[166] = 144'h0907f157dfd2018beebd1d19179509cbe5f3;
mem[167] = 144'he97a00151752e51e1a2dfc681950f1cff350;
mem[168] = 144'hf816e8d4e63705a20990e9f6ebe7edeef4c0;
mem[169] = 144'hf7aa19ea0ce7e0a102a1f1dbfe12e5a9e6f9;
mem[170] = 144'h006af01e0b95f27f18411bf816e40a0df9eb;
mem[171] = 144'h00b6e28df0a5e50916a20bd7fd061bb712a2;
mem[172] = 144'h08a3e2de1ff5ec02ed13f597fff8f1200b3b;
mem[173] = 144'he5e617580e39045c14b91a53e17ffc390560;
mem[174] = 144'h0145ff7ae560fb85e0a3fbf7f7380d0e0af4;
mem[175] = 144'hfec4eaf70ae9ea010378e16a0c571378e799;
mem[176] = 144'hffe0e6faff1ae942e22ce4331d3f16e30b74;
mem[177] = 144'hfd1ff2b81f07fa16f2b505540cabecd5fe11;
mem[178] = 144'h13fce1c6ebebe795fd7dfc54f89209c404cf;
mem[179] = 144'he225f380e6b41e50fc1719c11dc5e05bfbca;
mem[180] = 144'he310e57ff9bdfb07152c0797e754f68ee26b;
mem[181] = 144'h0a56eea6f24bf28c01c6eae4190d0b07f2bd;
mem[182] = 144'h0970e601dffb0049ebe0198a14321eec0982;
mem[183] = 144'hf2b7e5871e8bfee1037f1820fd15fcb9f62d;
mem[184] = 144'hfb39049ae5da11e01e3c0afcf690f239ef79;
mem[185] = 144'h0200124e1c6214dbe55d0a4b1605e45b1caf;
mem[186] = 144'h0532fc6e1088150f0ce31fb70644f1e6075c;
mem[187] = 144'h114f0be9fe55f7a3fae61b2a0c4e11ca09bb;
mem[188] = 144'he927086a1369fad415f309dcfc501adc1289;
mem[189] = 144'hf622168bf9b51d49f53a1daeeee016d41dfe;
mem[190] = 144'hf8dd1aca0f720d25f535ed6aebd8e3851993;
mem[191] = 144'h03d419901445f187ed1ce09d1e19e0470bf6;
mem[192] = 144'h0a0115bdf1c80085e9fefa65e46019041df1;
mem[193] = 144'h12651f66fc37e2a3ed5a0668f2951c8ded47;
mem[194] = 144'h14220a240960e652f7b40c4209a6f36cecd1;
mem[195] = 144'hf631fa06ec6807e90cd8e0f11506ebeee5f0;
mem[196] = 144'hef4201c903ed0840129ae16ce9adea35f24a;
mem[197] = 144'h09f7e8ee1e700288e979e147f8771117eb89;
mem[198] = 144'h1d5cf0a91b2f0496f066e808f7fffb19081b;
mem[199] = 144'h08c3eb4b0e2ee44215e9f64ceacce285eb54;
mem[200] = 144'h03efe69d0ceb0d80005c13b8043bf1e8ec1a;
mem[201] = 144'h0c821865e10eebf71e13016ae7c2117b0a13;
mem[202] = 144'h107418f6fe77066afb171ce8e024e3d70b36;
mem[203] = 144'h0317f12ffc8a0912e31b08aff63d0150e829;
mem[204] = 144'h11e5e4370d5b121206cafc5afbee124bf9f0;
mem[205] = 144'h02af1e9a01ed1121f4c3031c0e260bb7edf1;
mem[206] = 144'hec4c07b4e7180472e53718a11af30960ff42;
mem[207] = 144'he0b311acfe121bf110cef690f7b60f94fb25;
mem[208] = 144'h1a1ce3cef9f8e4f90cad11e70dfc1a6f1307;
mem[209] = 144'h19c00b5d0d74fc2c0f29e1afe350fb79f699;
mem[210] = 144'he5b9ea2ae83418fa14c5109a145006e015fb;
mem[211] = 144'h0355e676f73619190cf311ef140ff4bce8cd;
mem[212] = 144'he0e4167f06480632fc3ae2670e9817cc1b99;
mem[213] = 144'h04fb04c306730138074b0563fc8be7de15de;
mem[214] = 144'h00fe1513e200191ee5bffcacfee71539e938;
mem[215] = 144'hfcc109160e2afbd7f40de6dff80e1bfceb7e;
mem[216] = 144'hfe4914f2e7f41c8a19b508ffebcee641e136;
mem[217] = 144'h0f0be63df097e50807bde290e9aa17581817;
mem[218] = 144'h1217e4ea1c64f35c07d3fffa16d0f79c16dd;
mem[219] = 144'heeefeb2a14a6093c048402c5e93e1438fc2d;
mem[220] = 144'hf1f704d00960e72d11f20efcf2a81d05f669;
mem[221] = 144'hf5571448eae31e3fe99cf5b817b001cf0ef1;
mem[222] = 144'hfbcf08bf00a2ea5ffcd21c26e06eeae21fd0;
mem[223] = 144'hf3f60fe417730300f7781aa91be7e030e00b;
mem[224] = 144'hf018e640172e03f51ae6033efd0419d10557;
mem[225] = 144'h0a5e0bdf1c0af38d1f490d58e2baedac1673;
mem[226] = 144'h0ecd135fe534e2230267f990110bf1dafb1e;
mem[227] = 144'h03bdfe8517f81ec700a7ff0f1d20e336ef7c;
mem[228] = 144'hf86eed70e4cef2ed07f0e762eced13701331;
mem[229] = 144'hf266091aebf7fe9bf7ee132417d50df609e3;
mem[230] = 144'he0d21031025ff7fef141f36a11c8ec20ecef;
mem[231] = 144'h177b1b79033202f4014810f1f121e78f1203;
mem[232] = 144'hec991464088d10a502dafc31fdccf81bf108;
mem[233] = 144'h0922ee73fe87e5d2fcc90b580a88f6a41a62;
mem[234] = 144'hee53f4340b13e8e91c940855e093f0cd0f8a;
mem[235] = 144'hf7850d7cffc60d09e68c1779f74909c7e032;
mem[236] = 144'hf2f1ea6301cffa7ceabe009df4a313faf35e;
mem[237] = 144'h07b9e3280c89ef20f24618a0ef7ae1921c7a;
mem[238] = 144'hefe4057fed6e1195f464efd60052f77508e1;
mem[239] = 144'hf03f0bb8f5ff1e3002f6023919c41703049d;
mem[240] = 144'h07890f46fcefecc5023b0bcceee4ef460e11;
mem[241] = 144'hf61017b9ec7110080cace8eb1ef0f328e879;
mem[242] = 144'h19d9fa260a3115b314520451f7f2132c02dd;
mem[243] = 144'he447f2b706630968072ff8f9ebb8e940ee46;
mem[244] = 144'h1a0e14e9f90e120d1d2714660f3c0efcf530;
mem[245] = 144'h11c0eff0fda7052efc140b9f18a40bbc06e8;
mem[246] = 144'h1508f755ec191de2ec7ce820ee04f90a0a5f;
mem[247] = 144'h0c651581068716deec81195d1f1c01890b47;
mem[248] = 144'h15ed11b61e92eb2c146ff09cebbb0ec2f106;
mem[249] = 144'h11530997045c104a1a3ef17614500bd1e1da;
mem[250] = 144'hea151ad5fe7cf7cdfc71e1281397faeb1685;
mem[251] = 144'hf9b5f8f702c01fc7e9fcf6cd126f1ab60894;
mem[252] = 144'hf9470daff6cb11ade6990d7a1f2800b31437;
mem[253] = 144'hfcca1903f559f61bfa360ce0e87b0d85e2d5;
mem[254] = 144'hfcc21db4f613e3b01b120690170309a61386;
mem[255] = 144'h1569e6ea03d2f4e0e7351afaf0d6f932e8c5;
mem[256] = 144'hf267fa600ff3f451191a0333e7dc1be21d5c;
mem[257] = 144'h1eabf02feae9e0e7e3991b2ee319e5430d92;
mem[258] = 144'hfcf1f4f4e1c10077fd77ed28ec2712f401ca;
mem[259] = 144'h053fe10bf08513200fc414ad0ae80eae1789;
mem[260] = 144'hf36eed36f6b8f86f0a76f81f1780ff800f32;
mem[261] = 144'h016305c3e7edf9030655f30fed4ce228fe8f;
mem[262] = 144'h08170621ea59f686fa80f457e9ee03e7f4fd;
mem[263] = 144'h06a4f5b8e6c7f919e0d7ec13198812170288;
mem[264] = 144'h048b10fcf43e000017bf058805d6fa661a9c;
mem[265] = 144'hee5ffe2b10911b2f19fbf756140c06affd44;
mem[266] = 144'h0585f1b4eb67f85f1f79f7d1e0d1ecccff54;
mem[267] = 144'h1139f931ec3ce4aa019b0c311c8e18ae099d;
mem[268] = 144'hf44df80f0db8fc1a0236fde61fbd0e220163;
mem[269] = 144'h0de4f5fa142f16a91c441ee913a41cbcf88b;
mem[270] = 144'h1b3a067af50ce046033908a4f0de0f1be80d;
mem[271] = 144'h1512142b0b8fe1d3fe75ec970675e1610a32;
mem[272] = 144'heed618cf065d175de43316fef6451cb1f105;
mem[273] = 144'h03dde1b409f50e3f13421b25fc5bef4617e0;
mem[274] = 144'he4860fbf1f0de747e0e61c6309601d0febd8;
mem[275] = 144'hfe74189af6d7f9e8135017dd0f14fedb10c4;
mem[276] = 144'h1782fe6eefab1f06f10eeeaaed61f9b80451;
mem[277] = 144'hfe1ef7050c511ab5187b018e12ef1b810727;
mem[278] = 144'h06eef56b0b14ebc5e080f68cefcb1c86f123;
mem[279] = 144'hf8fae1850bd614ce1c740b1c084ff4a307b7;
mem[280] = 144'hf7e00fed042ef2661469f3ba11f6ef15febb;
mem[281] = 144'hfb980cc1efb2e6ede802132317cdec6afb1b;
mem[282] = 144'h013807eb0ab21d4715a3e09602ff1207e5af;
mem[283] = 144'hed3302df0912fdc911fd0a5ae52bfaadeac5;
mem[284] = 144'heef7edea1cedf8bd150cfca5e47a1044ecdc;
mem[285] = 144'h060ee4d6f4b2e430015c1cb70b48eef50f43;
mem[286] = 144'hf65b110be9c018c5f2ace2aeff21e1f21bb3;
mem[287] = 144'he1ab088e122aea57e9bbecb10526efecea57;
mem[288] = 144'hf4dae893f4f8ea65fb86f4680c7c1e87e664;
mem[289] = 144'hf5ec19480d75e92d1393f30e047ef312e7b0;
mem[290] = 144'hef710fc40284ff63e05200d2e03bfc70e53a;
mem[291] = 144'h0a5ded7618c9fedff58d1fe51474f5a3f60b;
mem[292] = 144'he96bf332e6eaed210e48f7900ea41735e107;
mem[293] = 144'he7e90e0e10830b4ae76deb260c400201f836;
mem[294] = 144'h0d2ffbd10ab7047fec4a16b01e8ae2c0fa3d;
mem[295] = 144'hfe33eeb714d6f08d022d0104f3dc079cf0cb;
mem[296] = 144'he61ff02df361173911f414ae09f0037b1fe5;
mem[297] = 144'hf1f5e97af9d50842f0761cc8fa510983ff34;
mem[298] = 144'h1641ff79fab61872ff3e02fdf96be885fb2b;
mem[299] = 144'hf08dff7c03b8e28a0fd2ea881991178b1b0a;
mem[300] = 144'hef211c3a1214e331025902c6fae00899f9a5;
mem[301] = 144'h09da1b3cf6b90396f4f1143710fce6fc1c15;
mem[302] = 144'h1fa6f370ec89e533e30e0575032f1c58f88c;
mem[303] = 144'hf7590ede0053fad01914eae8177407470ece;
mem[304] = 144'h022df33af855121ff42bed8ce9301f31eb50;
mem[305] = 144'h078ef992e1c612fffa0902cd075b01fa1dad;
mem[306] = 144'h0ed7eb22f7ed065deaa4f1aef21bfd3efdb4;
mem[307] = 144'h12500bc119a6e41c041aec8b0b96ef29f8a4;
mem[308] = 144'hf3d6f614e73011e703e9eb2c0740eb93fb3c;
mem[309] = 144'h15e1f588fee8f2f51ebf024d07b1ed071744;
mem[310] = 144'h023ff06b12af0ccaf105ebb4029de4231634;
mem[311] = 144'hf287094612dce384e65e171803cae4eaf427;
mem[312] = 144'hf8341430f5f50b2c1866f51de3d2e3e6e1e0;
mem[313] = 144'h14deed24e53715130695f900e777f5261a0c;
mem[314] = 144'h03b6006ae858ecfe1aa2fb0af277f5eaf038;
mem[315] = 144'h1a55053bf0330a2719f21e221355e6f4ea19;
mem[316] = 144'hf826e57f17abe5b60fa4e62302e1eab9ef40;
mem[317] = 144'h1d191713fa0d0b541d91fea1f3b3e20feaa0;
mem[318] = 144'h1202166af847f6bae2bd05f1e869ea7909ad;
mem[319] = 144'hffa4e284159ff3f900a6f78afc4be8c0057d;
mem[320] = 144'h0c0b17c11f290ee80278f9ac12931486f7db;
mem[321] = 144'hec55f42317770aa113b2ed77f60ae6f5e83c;
mem[322] = 144'he297e7860d3be5c6f76beeaa08df0663e1f4;
mem[323] = 144'hec29e9e1fca7136016b217a9f520fcdb0612;
mem[324] = 144'hfac41b63f11a16151e45119600d41b3ce1e1;
mem[325] = 144'he9f1fe900b921d4b16a2ed76f9e70477fea9;
mem[326] = 144'he3e8fb64009100420547e6320a881a07f32e;
mem[327] = 144'h1e5c02c5e65d1a75fcdef315118ce22c1625;
mem[328] = 144'he4cffaf607f10b9fe1ce03b80bfee6b31868;
mem[329] = 144'h0445f7e7eca8e552ebc51e62e1a6fb0619ae;
mem[330] = 144'hf06af5130bafe59eecc311db0147f41706e9;
mem[331] = 144'h0aa0fe7eeddb0cbfee18fef70f64e0be0546;
mem[332] = 144'he4dee6fb1fd3e599e93ae0f8f369f23df979;
mem[333] = 144'hf5f214281e48ff0c146b05a101dae821f5d7;
mem[334] = 144'h1832e112e5c0116c0f62f865f0c1e14fed25;
mem[335] = 144'h1f59e32b1363f40813bde9b61a46fc6fe0d4;
mem[336] = 144'hf85f092012d1fc8a0d44141d1064ef24176f;
mem[337] = 144'h0bef0d2cf4a9fdb71ac010e51a3efe01f2bb;
mem[338] = 144'hfb2beb231ca21e9b0df71cfd05e515eefbd7;
mem[339] = 144'h1d891e5bf135f67805b4f3aee238ebde023f;
mem[340] = 144'hed74e1edf10dfd86f341f51f1d66149c1230;
mem[341] = 144'h1111ee530df4e10cfc420bcde9590c1efd81;
mem[342] = 144'h038fe24712ec0d38e76fe1210b140c6a109e;
mem[343] = 144'he532f1fa1a970d5b0fe8f369e542e4c4e3c8;
mem[344] = 144'hec5517a2175ae76c1edb1a080a5cf808fe23;
mem[345] = 144'h11c6f54918ede141f101e65ee8fa13ce0845;
mem[346] = 144'h0186e0fd03dafd51ff2a113cfce1184016f4;
mem[347] = 144'h111ee82910a2e73ff96eef72f2260d0f0ba0;
mem[348] = 144'h133c17f719f2eb3ae95605f8f0c7f9330dfa;
mem[349] = 144'h1c8ff0faece509cf1d0eee8904b01df2058d;
mem[350] = 144'h065916e70597e4e4f6c1199bf5a00709e7bf;
mem[351] = 144'he6c719f818b2e5241c6c1bb4ed171282f7ee;
mem[352] = 144'h103011eefb851df0f62a08eb005bf7edf10b;
mem[353] = 144'h0fb7151d0c1df936fd1a08beeb8c086014c3;
mem[354] = 144'h02930827f87709cbea340c1ff4d2e1ff03b4;
mem[355] = 144'h023e002c0372165b0087fa52e7b1f4c1f559;
mem[356] = 144'h111e0e151be90b77ffcff436ebce0bf11ec6;
mem[357] = 144'he313fb2aed9fee921553f8dbe2faf0eff364;
mem[358] = 144'he448e4fd056d1accea321312074616a30320;
mem[359] = 144'hfb69f75af7430bca0218ee2d0e9b1690f5dc;
mem[360] = 144'h1c9be944ee540728183ce3aee3691cefea4e;
mem[361] = 144'hf9c6f6430a2519daeb441b160b580d771797;
mem[362] = 144'hf04c076f1963e7d2067ae97d1a2203190d2d;
mem[363] = 144'he9301434e07e055ae90dff620c44e62719e1;
mem[364] = 144'hee9310ab0256075d1b72105ff6810f3afaa3;
mem[365] = 144'h0ff01119e6b3ed33fa95fcad131f0118f422;
mem[366] = 144'he6851739ed6eff7df1700bb707560039f04a;
mem[367] = 144'h1c5afd63ec381e2603a7021affd914d31299;
mem[368] = 144'h1d2403331604e097e04bf8031a091a4104bb;
mem[369] = 144'h1feafd1bffc4110a09ed02ebf37816e815fd;
mem[370] = 144'h1d0c15e20c59fd83f1d70d4e1f4bebfc08e2;
mem[371] = 144'h1a87190deb721f7a169f143ff228f0e516b3;
mem[372] = 144'hef86f814ebea1305f22c0e60ecd9fe070c28;
mem[373] = 144'h10df07c9e8d714f0f2d0eeb0efb9fbc8036f;
mem[374] = 144'h1021f58300e21815fb2ef075e44411611166;
mem[375] = 144'he537062af4c310a41b67e8f3fcf713ca1c4f;
mem[376] = 144'h13b11cdef859f73809880b7b10dae59c09b6;
mem[377] = 144'h0be0072d0897fedc00a3e03e15d9f3390ab1;
mem[378] = 144'he8ff1eeaf0d913a103aee9a0e303e3a109ae;
mem[379] = 144'h013fe1fce9031ad9eead178ee632188a0afd;
mem[380] = 144'hec56e60a1bdb0a1609b3eace10d705230779;
mem[381] = 144'h1a9eeb610c7aebf0e891032616d105cf179e;
mem[382] = 144'h1b4bfed11bc8f7a5188b15ef1441f4ffe899;
mem[383] = 144'hf156f65de4ba00e0131b012ee33bfc9df968;
mem[384] = 144'h159bf6d0f59905b0e7f8f5d1f5fee215e6e3;
mem[385] = 144'hebc80a0d12dce7acf21819b00eaf0fd31232;
mem[386] = 144'hed5f00a50688174809470a0be7e31c64e231;
mem[387] = 144'h09530e7f1706ff080bd4f79715a61521f0f9;
mem[388] = 144'h18b705a2007aef14e4c005700a2f18d411e7;
mem[389] = 144'hf66fe5d9fe7211de011504c6eb12120904d0;
mem[390] = 144'he248ed1af8b2f1ade3a5f6c4fd811cec116e;
mem[391] = 144'h169e154d1d50e210f93d1d62e947f45fe8a0;
mem[392] = 144'he7fee9dcedfbfa380d5e0d59e23819e0f6c9;
mem[393] = 144'h152f0083e0f31438088c146c06b7e689f692;
mem[394] = 144'he1eb06960540e93917df0255f6bd14041244;
mem[395] = 144'heeceef41e29d1c35f7af14121ed511c70401;
mem[396] = 144'hf0a7064d1911e8f518efed48eb8ae29eecd8;
mem[397] = 144'hee20027ae2c417b2ffb408480d480e96040a;
mem[398] = 144'hf25e0ced160c11980fcd17bafbbc1866e9ad;
mem[399] = 144'hf868f0dc02a1ecd918f1f8720e7c17affce6;
mem[400] = 144'h1405002ce598f8f3fe0cee6810e3ed4df5a6;
mem[401] = 144'he1e3f77d1a47f8f6e1cc12bce4dcea8806a3;
mem[402] = 144'he772ea9c119ef0d2f26211da0f191cab0d6f;
mem[403] = 144'he9d2ffd1eecaf6cfe6c8fb3a19b00c911bc5;
mem[404] = 144'hf30bf51ee9721024e72111c70f4d1edf0645;
mem[405] = 144'hfd6fe98b2001f3a10fb9e833f0a61b16e92e;
mem[406] = 144'h1d530eff04ce1b82fdc912fff674f8371c45;
mem[407] = 144'h18920df7e63f07d1ea140b89e59f0e331067;
mem[408] = 144'h1dc1e271fc8bec8b1c3c1c90196affe8e63a;
mem[409] = 144'h13e2f05aebf31b87fa4017d2eadcf668ee45;
mem[410] = 144'h0c3f00b704aaeec70f8003efed5d0a2dfa9e;
mem[411] = 144'hf7c2efe50afbfcf1ef12f45319870baee16d;
mem[412] = 144'he50e0d4c04890d79019f1955e000e2c7e2a0;
mem[413] = 144'h085f156b059fe152f5f501eee3d9019b1e61;
mem[414] = 144'hf35c1183eb6a15a71c230091e1191e0efec6;
mem[415] = 144'h09c2e8c70cc6eeabfa3d031d1222ed1df65b;
mem[416] = 144'h17e8fc590bc41cacf8780f1a0751f3e7e3e0;
mem[417] = 144'heec01fca1123ede41d440a08e54ae2270691;
mem[418] = 144'h095c0db705e114bcf49b0526ea06fcfeead6;
mem[419] = 144'he35706ddeac2e37b0020e5d6fcccf559f8f3;
mem[420] = 144'hec34175b1aed1ae2e4d2f703f7f6e212f237;
mem[421] = 144'he31be992185f175af857f23b1d3af9380e29;
mem[422] = 144'hf7edffe3ff8cec1f1cdf043d06bcfaf3e735;
mem[423] = 144'hee7be877103f0112162d138219681649e443;
mem[424] = 144'h0698f8c7ff9f1528fba71d430d43f04bf6c9;
mem[425] = 144'h15f61f8de198e8dae60211d50458174eeaf2;
mem[426] = 144'h04a5ff9de44a0d3ff4cff3faec06e780e732;
mem[427] = 144'h1bda196bf16c1f1b05001bed161ffaf710a2;
mem[428] = 144'h1024feb002531e69f9fd02faff56e7a003a1;
mem[429] = 144'h1783ebe8ed2deeb8e35902e0f2121cafeeda;
mem[430] = 144'hfc15e4500adc024dfaa8e5dcebe1e537fddc;
mem[431] = 144'hea591190e0f00ac3e679fd7deb1ae9061aeb;
mem[432] = 144'h0ae601d6e0c9eeb9eb4fe13a0b5512a309e1;
mem[433] = 144'he724ec92e59a0c6f1056e43c0e94f62bf2fc;
mem[434] = 144'he6f01a0df813f50ee9f20035fbd113e505fa;
mem[435] = 144'he0f7f65be1b61a7ee1320ab81f4405220bb7;
mem[436] = 144'h0e5816b81b7c1fa81fc2ebd31e7814c90fc3;
mem[437] = 144'hf2c5e5aee27e1b59f0fbe4e306f9f8f6ecce;
mem[438] = 144'h1fcbe46003aeeef318d5120d072df0aa1758;
mem[439] = 144'hfea6ee50f80b048bea7b0251fd0fe3f21cac;
mem[440] = 144'h0b4df27e10cc1c611a4b1436e5b8f3100a5e;
mem[441] = 144'hf64c022812dbe91af65919f816111857e040;
mem[442] = 144'h01e5ed700b4411d7e2c9ed18ed29f1e21356;
mem[443] = 144'h0647fff3093a15ca01f60910098b1d02f91c;
mem[444] = 144'hee2d19ff01c0e9c114e813a4f1ea1863e37f;
mem[445] = 144'h1bf41f0c018c118b10c60237f5a5f8601687;
mem[446] = 144'h1919eb871c87e2dae62610da0b59e1220f09;
mem[447] = 144'he6ff13e3fd010959f630e3440f27e72a0d88;
mem[448] = 144'he5da09a1095efc3214c1e71c03d7f5060491;
mem[449] = 144'h059b0987f533efa60766ff03eef114011b52;
mem[450] = 144'h1ef2edfd16711c3ef8cf183d15431b7306eb;
mem[451] = 144'hec9101adf4a30d1efc530ecde22af26cf19a;
mem[452] = 144'h1d3c0314e8c01882066004b7e2410a320c68;
mem[453] = 144'h0fb40b641cb40feaf0c9f8ea06f30aa1f1de;
mem[454] = 144'h108ff8f0163e01e319e3ff34f378ffc7160e;
mem[455] = 144'h08dfeddfe5ac051a16a8149318e10a7109b6;
mem[456] = 144'hef88f5c0e9c519a91ee61749f55d06b8e959;
mem[457] = 144'h1c15f406f34717da01d3f68ef8cf1ebfff3e;
mem[458] = 144'hec7208dee0790c0bf6af07a2e75d01f7f608;
mem[459] = 144'hea37f691eaeff8e2f55300d70bc2ff34fcb5;
mem[460] = 144'h07c9e5db0d45e5f2f288fdeafa9cee66fb92;
mem[461] = 144'hf9f815791000fc95ff66f0a3ed820422fa32;
mem[462] = 144'h0505ff2fe4f7efd2f98404620c3a1b01054a;
mem[463] = 144'h1cb9ed03efa61fef0f59f44ff3510723066a;
mem[464] = 144'he1d31b67f7001ada14aff091f0770c38ff28;
mem[465] = 144'hf059e391fc1813311918ef44f9b11e131693;
mem[466] = 144'hefe517beee73efa01954f926f7090b0e116f;
mem[467] = 144'h01c613010388fc0d1a13f3411701f0e6e1ca;
mem[468] = 144'h19b2e2c717c80038127efeebf502fcb1fc52;
mem[469] = 144'h1b4403641900fc3e054b17b6f00a1d190c98;
mem[470] = 144'he556f05d0b93e852edbdfc2115b4e081f206;
mem[471] = 144'hf9fef0681ea7ed6c15f0f0cbf9f0149be6a1;
mem[472] = 144'h1bd50a1a18c5067ffc28eabbe8d8e9080ea0;
mem[473] = 144'he4a6f9e3ff0ef3c71f8d179f0750fbc9fea7;
mem[474] = 144'hfd010f3704eae79410a1fdb3f64a0ede0cff;
mem[475] = 144'hfce11ac7f18b1858eec7e8e4fd8e125eee9f;
mem[476] = 144'he55bf32de06dee91eac7e2f118e2191afb22;
mem[477] = 144'he3990299f8e40187eabdeabb10d9e649f6b3;
mem[478] = 144'hf37816b20506e87be6e60103e984f10ef4ef;
mem[479] = 144'h12c818e1170907cafb4af688f45af6f81755;
mem[480] = 144'h1348e024f4c6113ce9f4071d1d69fd54ede8;
mem[481] = 144'he670f3a407e1f37de52f00e21a43fff810d7;
mem[482] = 144'h06ceed8e13011d4118d1ef87e4e1f7d4e39a;
mem[483] = 144'he973f18314c41de8e2d1f59f01d4f0a01c2f;
mem[484] = 144'h0cd60226e0cae060171ffafc09a904b8fad3;
mem[485] = 144'h102b1395ed940255fcb2072f123d1ab8ebec;
mem[486] = 144'h00ce107ee2aeed89081af5ffeb0e1823ee66;
mem[487] = 144'he5d519120b4b14fcff160c900345e6a4f98a;
mem[488] = 144'h0222f7ce1d80fad3f03df4f5ef3de788ff99;
mem[489] = 144'hec431281ff7ceab3e6f7072d00b2ebf6f166;
mem[490] = 144'hed67f01710ce0aa91dde076107db14e1098d;
mem[491] = 144'hf471ff6fe1870683fc3407fc1527fe821319;
mem[492] = 144'h12850638e0dae5a9fdce0365e05e122f013a;
mem[493] = 144'h130b13b10df41069f5450edf0e67080e041a;
mem[494] = 144'he1bb1dfae9470874fdf01d1d02acf506fb18;
mem[495] = 144'h1626f641f34ef9f812caff6116dc08df0f82;
mem[496] = 144'hff86fa86fb3bfcdc0aece41d1d021cdb034a;
mem[497] = 144'h0640f757f32916f6194f0e77e392f91de05e;
mem[498] = 144'h1445158c1fcd00b1f931f20603a5f9f716b4;
mem[499] = 144'he4aef2bb13790e521c7d0eff1e6e0b55022c;
mem[500] = 144'h141014d10e36e0f714eff44fe2851311e9a6;
mem[501] = 144'he94bf99a1ed81801fc93f779e0b9f794fb00;
mem[502] = 144'h177c183e1985f013e117e384e05af513fe6b;
mem[503] = 144'h0ce40f0d150bf46011881677e588e600047e;
mem[504] = 144'he0900ffb1c8ae081084b117a1e26e76efe02;
mem[505] = 144'h0328e15de3da15d2085d1ff9fb03f7c21112;
mem[506] = 144'hfe8c09e7f6810118115be065ed61eeafe00b;
mem[507] = 144'hf659000e198ee2d5e4a1e7c007affa741a85;
mem[508] = 144'he1341dfe0f770d4606f70843169b0f1be516;
mem[509] = 144'h1b0ef7ccf146096c13690993fc3df78ff72a;
mem[510] = 144'h17191b341fce04100d490f32e5b2083fe29d;
mem[511] = 144'he53be4e2e3a01ad3e0a205c2ecbce213ffcf;
mem[512] = 144'h1d9b0fd4efda1bfde5f0e44beec912d5e176;
mem[513] = 144'h0e69fd4be53a0d4016991df7ef370060e029;
mem[514] = 144'h151f16fef20104220b3a19e8f188fc15f898;
mem[515] = 144'h0382f646e18f09feeb781f0e182401440af8;
mem[516] = 144'h1773043e183be6241bf71e3fe8ae087f0294;
mem[517] = 144'hf63504c1f0b11e921e47097ce7e70404ed2e;
mem[518] = 144'h0a2817acf0f1f33d11aa0c8feddbec5cec4a;
mem[519] = 144'h122900dd1da4fc671635e59011ba064e085f;
mem[520] = 144'h1e160f8cf941e3150634e2311e0fe2230465;
mem[521] = 144'hfe44e7b90de8fdc60679f1cfe665f8a9103b;
mem[522] = 144'h0e5e061014dee331f248fefcfc351b0af0c0;
mem[523] = 144'h115dff5ce47bf9e0fcb51601186ce7ec0d64;
mem[524] = 144'he91f1049fa891e26e16605a7f6efe50a1504;
mem[525] = 144'h0292fbbfe8d30f61ead01244e7b20d6e0a0a;
mem[526] = 144'h1bb612bc1eebf88f1f6afa95ffa41068f204;
mem[527] = 144'h060ee1afe29d1cbce1ea18451e660487f826;
mem[528] = 144'hf57113b11510f29be160fc0c00beee231b8c;
mem[529] = 144'h0728e82a178214b305fae431e7730ddd178f;
mem[530] = 144'hff4c017f0d771f99f0240cf9e8730b6ff993;
mem[531] = 144'h1ecd180ff7c600f1f7a60cb7ea53e4e906e1;
mem[532] = 144'h18d8ee08f8cc125ee24bf087ef47128aec91;
mem[533] = 144'h1933f1620833061c12df078109301339e8de;
mem[534] = 144'he467edad03b1e86be0c5e146023bf2251aa8;
mem[535] = 144'h0bd8fdcd0868ebcef99f1dd4e836094af154;
mem[536] = 144'h1854f54511ef0138e0ade27613a3e3ce0901;
mem[537] = 144'he4ddf276e012024511baf2d911a6ecd1f328;
mem[538] = 144'he27d027f13611a2bf734f603f3e9f784eeeb;
mem[539] = 144'h0bf30b96e5ae145607bc035be403f9f71f72;
mem[540] = 144'h03de0c84090df9411963f2c101acfa83f17b;
mem[541] = 144'h15b80dcbec590ab50563ec820cca0de8f478;
mem[542] = 144'h0505f9251709f1be11111b01f85f071bf37a;
mem[543] = 144'he379e10bea6a09d30528f5171b33136317b4;
mem[544] = 144'h1984fb0f0f7bedbf112c1fc9ffa0163ce471;
mem[545] = 144'h0c89164a0efee7490f31167912481b35e536;
mem[546] = 144'h10b0fe8d0a8a11581ccd16980cc7fdc4f4d4;
mem[547] = 144'hea6ce5f9ff7b1822ed23e5c1f69ee393100e;
mem[548] = 144'heec0f4b2efc6036ee8f1044b1700e3d00ff3;
mem[549] = 144'he91306d1012f0589ed7ff59c19b2197e1415;
mem[550] = 144'h1b36fc7b071dea75105ffaf7f5eb1ccef435;
mem[551] = 144'h0cc4e1cfe1d1f0e703d50cdce753e48b0f5e;
mem[552] = 144'h096e111b15a1fecd02521fc21b141190f10d;
mem[553] = 144'he1c519ba0dee1f1ffdf4177bf0b61548fef4;
mem[554] = 144'h0838e58ce6b319140f12e7dd1984e26f14fe;
mem[555] = 144'hee31eea60094f513ebce10910a11078cea85;
mem[556] = 144'heccbef53fa10fc58e6f4ef4e1490127cff93;
mem[557] = 144'hf2bde9f4f22afa90e265f9281e5ce3c3e8ae;
mem[558] = 144'hf601eb06fc9dff2ff87107a50cbd13c9e45a;
mem[559] = 144'hfd25e38d1c910df2f7a1070eea40fb3b1060;
mem[560] = 144'he2150fd5f0fffe711d42fc8d0197166d1146;
mem[561] = 144'h01601bf6e1890819f7a6e73d0ff4e4110f55;
mem[562] = 144'h1a9118f4fa8df41507fbf83cff191d02038c;
mem[563] = 144'hea06ed3bfdd4e3dae61efe21e3b6f08f1ece;
mem[564] = 144'h0818e42ae7260e0d0e6ef6881a87f8ec0dcd;
mem[565] = 144'h167a1a70ffac18831cb5ea99f8a81b28f506;
mem[566] = 144'he285e1741480f15cf535186dea9c0914e6fa;
mem[567] = 144'hf52bfb32ffbae4b2011be4d6042b1d3bf7ec;
mem[568] = 144'he5b6f13210cee0d1013dee180baa0e6dffb5;
mem[569] = 144'he34e0073fd7de723e95af540e393f695f98d;
mem[570] = 144'h127a1f4ce41ae779ee68feb71772098800ca;
mem[571] = 144'h1e6305c7ea50fdc61d6e0e171dca066d0f45;
mem[572] = 144'h0b2afb541fda141ffcb1fde51c72024be67f;
mem[573] = 144'h1d880282e779e782f95ceeb0f4a719301881;
mem[574] = 144'hef75f401fe6d050bec3403810f201f41fe50;
mem[575] = 144'h1621eff0fff9123e1565125d0c9214e6f3df;
mem[576] = 144'h0af8092b01870afcfc20ec1a16f215561ec7;
mem[577] = 144'h0925044a10a7eee3e2fa099ff6abf7ef0cb1;
mem[578] = 144'h19aae42affe4e3b4ed3f0883ebb2f6b4f2e8;
mem[579] = 144'hea7af361e2acfe2dfbb308aafc6cfc280e92;
mem[580] = 144'hef9df7ed1632ee9f17d0f3f8e07dfae50d16;
mem[581] = 144'hfe900499efc91295e3ad1c7b111cfa70fec1;
mem[582] = 144'h1f6811b7031df5c7e669e01b0729f1e3fc01;
mem[583] = 144'h0b17f0c1ebc20ff9f2b21c581df7e7421177;
mem[584] = 144'h0916ec66f8ecfd771afa0aaa093919831720;
mem[585] = 144'hf93c1a4b0d0208b5ede2ed65f732fbabf83b;
mem[586] = 144'h1df0e501ed46fb2e1a00fbf0e4db1457f820;
mem[587] = 144'hecfa01e6ed491d5dfb78e998e5681a70eb3d;
mem[588] = 144'hf0080571fb111d0aea52f9c5e96a1987f807;
mem[589] = 144'hf41903efe3dcf412f6871e4d12b61ba1e6da;
mem[590] = 144'hea77e8c4fbc8f970fa80e478f6f1e811f2f2;
mem[591] = 144'hec780134153cf0f1ffcd1864f2acf60d0aa2;
mem[592] = 144'hfd441b6f0c6d1e08f63ee7260bc1053c0fde;
mem[593] = 144'h0907f1f70873e432f28af9b31a820e18ed38;
mem[594] = 144'hedb6009b1cbfe2d2e705e205e67bf5b3f76f;
mem[595] = 144'he506f6800794f3f2f1cf01a5fc3bf23716f9;
mem[596] = 144'hfc56f08c0a38e0d0f7f1e09aefc20a810f20;
mem[597] = 144'h1b441f1de46800f7e15300ff18d8ed06e41e;
mem[598] = 144'h0ccffa3de19fedb41a480086f246f49602aa;
mem[599] = 144'h148ff77507a7f96d1aff1d99fb37e0540f80;
mem[600] = 144'he4d9e295f654e247eb1efd40fff9ec750c55;
mem[601] = 144'h1e3ff17c12b1e87d17b1fde0ed2af5ae0070;
mem[602] = 144'he0d6e5aef0dd06cbe1120b64fa65faf50963;
mem[603] = 144'hfc12033d063de95f190809f4ea7d1391f12d;
mem[604] = 144'hfa71fcbae63215a5160c1ae81d99e0b9eea1;
mem[605] = 144'he9ff01700e50e8c2e6021ec5e5e01716125f;
mem[606] = 144'h09e4029a1aaef89d091315121eb6ee36fe59;
mem[607] = 144'he36d169cfd4f01291e78f43d1f55e4af0508;
mem[608] = 144'h0734153ef2260b81e63bf183fb2701faf406;
mem[609] = 144'he12ff5f608181aa0f6b5e9b91d5afb050e34;
mem[610] = 144'h030307bb1d01140704371ae2ece71955f656;
mem[611] = 144'h0dfa0e8204faec71e671e909f4e90b6d1f60;
mem[612] = 144'h1219f0ae11e6e7b2edd60ac30706089b0a07;
mem[613] = 144'h02a6e123ea8f0381edbb1cd7e4dceccde546;
mem[614] = 144'h1724077415cce4e411d00febf354fb83e301;
mem[615] = 144'h1897ead5f7ea07b8f9ecf8e5ffe8086e1cd4;
mem[616] = 144'hf32bf9531e7e10fb0689f1721f35f3cc015f;
mem[617] = 144'hf6e81556e0751a091c8805b20bc1e9851127;
mem[618] = 144'h19fbe0f9ff40f85311f70a5c1a1e1382ea59;
mem[619] = 144'hfd9800e2e033e0960e3003130991f534f0c1;
mem[620] = 144'h06e9f656031af2690666e1ed14c3f8b6ff08;
mem[621] = 144'hec341e3d200e0d08e5eb1fa30970eb9a0675;
mem[622] = 144'hedadf633e2cbe695e4f0e3ffec9f078beaf8;
mem[623] = 144'h1151064311c21028f9a8e4d5ec2afd4217fe;
mem[624] = 144'h0950024a17c3192707b8e064fb37e4770f28;
mem[625] = 144'h0e5f06bc0e791672185d11581250f7ccfa7b;
mem[626] = 144'h12390ef30ee8fa5ff18ffe11e8a002e90856;
mem[627] = 144'hfc9018baf322e9b5fffef1a91a861cc71098;
mem[628] = 144'h0dd0fe3df6f3088304dd18af1f0218a91908;
mem[629] = 144'h01cdfd540a1708fff319fe0ff691e043f4b1;
mem[630] = 144'head41e411d34188ae8c90b26001019050353;
mem[631] = 144'h12160e9d081de9081a3204f21258168de670;
mem[632] = 144'h080d0f52131bfb7ee084f2d20e6ceefb1111;
mem[633] = 144'h01e80797efb31aede711e0a4e7d2eedef931;
mem[634] = 144'h1b281d151126f0230836e881e5d1ed3e04f6;
mem[635] = 144'he45e07af0c0508831fd5e2d7ef7c05b3e271;
mem[636] = 144'heeba15a0f6c914c2f5be0f6606cee755ff02;
mem[637] = 144'he82bedeaf1550c1200f8090f1a61f44d1b75;
mem[638] = 144'hf82b1e0fe73003a2e2ddfb85ee6cf1d7122c;
mem[639] = 144'hf3b7fe76ed9c15f902d2f09ef87fe4a510e0;
mem[640] = 144'h0a06eeca13bb0448f862f0241aef16d0f64d;
mem[641] = 144'hf634f9b40659157eed421671f2ffea42fa71;
mem[642] = 144'hec72eeb8f89ff896e48e0146f4b90ff40a86;
mem[643] = 144'h00a6e352fbdb19abef491f26ffa71187e950;
mem[644] = 144'hefa8e611ebc9e0f9e1a4faf71ead0723ff6e;
mem[645] = 144'h15e5003e0d01f4d3f7af1b6d1db21ef2f44c;
mem[646] = 144'h0c30f83814a3e9211d67eb4f01d4f4af05aa;
mem[647] = 144'hfdd6f41415d5f780fef0144d0560fc7ff45b;
mem[648] = 144'he1d40e85e4351ce613cb1b9ff84ee0c6e630;
mem[649] = 144'h1042056ee5c60358002fe629ffc407c3092f;
mem[650] = 144'heff403141f58118efe77ee701b6ef3e80475;
mem[651] = 144'h1dd50c51fc52169c18e1f133103b0ac3f89d;
mem[652] = 144'h02951576f2ce1f93f2710a1df51e0e72fe32;
mem[653] = 144'h199decd31a39e249f35e1243e4adfb1514cb;
mem[654] = 144'h0d661359ec93f3e2e13c15841309fa3c1fb2;
mem[655] = 144'h0f050532e8dce2230d3ce7e413f1fa08f30a;
mem[656] = 144'he70ff07b0bdefe2ee40ae5f0e32b1ed01659;
mem[657] = 144'h0f05f8fc1e75e471f54ff188085f08bc163b;
mem[658] = 144'h0fcde166e291017bea24110b1cd6e7fe1f7f;
mem[659] = 144'h06bbe507e8bfe486f66112df0d7508b7f4e2;
mem[660] = 144'h0f39e40be0a71c2de2c916f307a10762f5e0;
mem[661] = 144'heb7f0db116b9f553164c128503e31ae9f596;
mem[662] = 144'h164b0c13f98f1368f5601f44e0e8f76ef1a2;
mem[663] = 144'h126e09eb1026e98ffa2de4e2fe0917eae007;
mem[664] = 144'hea12fefc0a7d0465056c1754e506e6d8fdc4;
mem[665] = 144'hf71c07b9121cf503f3660e2009d411e1f398;
mem[666] = 144'h1dd906c8f6961de7e010e893184617d9fc0a;
mem[667] = 144'h1515183de73006b1f13502b1f208e4c0e0f4;
mem[668] = 144'heace1b6410490f04005a0c50102c17f51d09;
mem[669] = 144'head2ec01e37417e20859e23df9dff98be023;
mem[670] = 144'h0479085b1983e7d61639f598f72b05c4080d;
mem[671] = 144'he69d1fb7f787137105a31efdf5461ae5fd00;
mem[672] = 144'h1c34e217e6d7efdaffff122117bde42e100c;
mem[673] = 144'hf88afcf11663ed370369e43cf139f45def28;
mem[674] = 144'hfe70e8e5054f1919e32bf585020efd021c70;
mem[675] = 144'h1884e0edf32f1d5603bb1bbc0a89103be1d8;
mem[676] = 144'h1a1a1441e5801ff91bbe1cac1cb118231d9d;
mem[677] = 144'hf1ad0c33f145e9801c46ffa2165f11ac09dc;
mem[678] = 144'heeb0fcf300341c9506f3190ee78f11a1fac8;
mem[679] = 144'hf18b0a6bf808f6c80cbe1761fe47146effde;
mem[680] = 144'h0ea1e85f12da17e2f21fe6430ee3096f0f8b;
mem[681] = 144'hedcdf701e1061a7011aae33a0202eee6fa67;
mem[682] = 144'h0133e0d1f8740261e4b40259f330058df118;
mem[683] = 144'hf11df9f31b77ee98f34bf094fa380573f647;
mem[684] = 144'hfd5fffdcf690ed21fed5e2d217331da9119d;
mem[685] = 144'hf781f73e116909a4eb3ef45e161ce6690a3c;
mem[686] = 144'h071ce0c1e6541e1deb9dec30eaa5ebb4e7a8;
mem[687] = 144'heaf6e69207c6e1f000b90a46f7f9f8aff094;
mem[688] = 144'h1fc513d3fbcef166122d1d39f4e1eaf2fad9;
mem[689] = 144'hfaa10ba11714f601f41815a8eaabf506ec6e;
mem[690] = 144'h0554113f0424f9fb0b930810efdae4c8f66c;
mem[691] = 144'he7cdec5f10b70cc70305f648153c0fca0c71;
mem[692] = 144'h15e7e461f516f835f9b5f812f7eb1114e7ff;
mem[693] = 144'hea011f7de0fb0e25e403e0cc168312d1faa5;
mem[694] = 144'he7fbfbd50903f53b04350c6ce8e4097bff27;
mem[695] = 144'he44c019d0bc0feaf15c2eb9bf5afeb251da9;
mem[696] = 144'h02040bb90f33043ceeade88700d1f6db1942;
mem[697] = 144'he0e9fe34150dfb6d0e80f4cf1d17e15ce77d;
mem[698] = 144'hef6a03231e2611b5fd58e359e05f101b0c42;
mem[699] = 144'h1a4d06a404761da41172fd9afe7fff19003a;
mem[700] = 144'hf0c40cc7e6550dd416e0ef38fd41f310e9c3;
mem[701] = 144'h0fd3fe99109d1decf7ece5a9fe22f140eccc;
mem[702] = 144'hf793f970ea38146ff5d61676fe9f1790f495;
mem[703] = 144'he115ef400f75020b1c650f45feb8e2be1fd3;
mem[704] = 144'h09830b93098e0349f5ae0c2ee6a00ddfe307;
mem[705] = 144'hf27bedc81facf2dc1062078201b9e8120d63;
mem[706] = 144'hf0ad1e11f6bb06ae1208f4ecfbfc0a74ec5a;
mem[707] = 144'hf294e1afe240e0c2faeded5ef08405811d5b;
mem[708] = 144'h1e2cf30cf341194b123ced03ee901001ed5a;
mem[709] = 144'h122ff13403b0f790fa23ef4b0e54034e153f;
mem[710] = 144'he346ef850bf8e32b1e88e66510c6e05306d0;
mem[711] = 144'h1f000484e3570433ec36156b082ee742e17f;
mem[712] = 144'hec96f0d8ffd8fe31e6150b0b016e16cee63a;
mem[713] = 144'h0afef418e459120ff10af2e00d8805a70ddd;
mem[714] = 144'hee440060fdabe8b605e6f05e1fc510521e67;
mem[715] = 144'h0aaeef72f16008330bf0ff6de11dee3801fe;
mem[716] = 144'hf166ef09f4eaeaeff3a21851fe71e13e024d;
mem[717] = 144'hf372060e07aaed59149906871b42f7eb17f4;
mem[718] = 144'he5c30fdcf58f13481bbbe407fe5d1eb51503;
mem[719] = 144'h1fa713eae2f6f4580943ee27e09b0a5de6c9;
mem[720] = 144'hfbacf2a4f0a5e1e8f121e70f10be0402ed6b;
mem[721] = 144'hf81af5e218d6063f1ccb01d7f350f0b013fb;
mem[722] = 144'he56ef8c11855e61113acf3e90ad20d091adb;
mem[723] = 144'he3fefe01f14fe056f8b80b9b113b117d0eb1;
mem[724] = 144'he9251268006c05c3ef87eb78045de767e9eb;
mem[725] = 144'h0745034fecfb06e51c9bfc691c8b0d9317f5;
mem[726] = 144'h08f5eb3a12901b491ff31858ed45e63115c0;
mem[727] = 144'hfdd211a713a804c1177d15d3e814fd280023;
mem[728] = 144'h1ae1f79c10e20684022efab31430fefff3a6;
mem[729] = 144'hebc8e478ec5eeee3115a1b3e1668ea1a019c;
mem[730] = 144'hfd011367ffd5f3f5fab5fc870543e1cd1a00;
mem[731] = 144'heaae0088e09aecb8e8f409dd0c571a7df9fa;
mem[732] = 144'h067ce2e811dff2431ef7ef8ae24ae1500e4b;
mem[733] = 144'hfdb01a4809c9eeef0213fa6d0c621fe1f3bf;
mem[734] = 144'h1c1eff7bfda0e350f144f706ea301e401dc9;
mem[735] = 144'h1a0b0eb31bdef2e3edc401f607a4fefaf955;
mem[736] = 144'he211004014bfed70e0eb1925ed5e0ef01611;
mem[737] = 144'h0aa60ca80b271e071cf8efa100391af00cec;
mem[738] = 144'hf3151f9407f8f581f0f70959030d1ad0f27a;
mem[739] = 144'he930ef941fc3169cf85cf6bffa47f91f0f27;
mem[740] = 144'h16d8fd35f8be157206f2f39a03d8ed1013b0;
mem[741] = 144'h0863e3c71ad1e069ee4118d30c96e402032e;
mem[742] = 144'he501093618241193fcef1a21003aefe71953;
mem[743] = 144'he98f1bfe0e5c13280779008d03b11bb0faa5;
mem[744] = 144'hedc71ddb040e1bcde8ce00a7156aea02e806;
mem[745] = 144'h0252ef86e4e1efd215d60ce1fdbbe87ff8be;
mem[746] = 144'h1e190096ea75ed920cf4ecf1f19f091b0b16;
mem[747] = 144'h123716ccf6160b81f284f77e0486e1ade93c;
mem[748] = 144'h0f9bef65e645ec86021415071700e7c8e578;
mem[749] = 144'he384e56e0ee8076df0170b6eec9afb57e648;
mem[750] = 144'h159c0fc70c69fe31134e02a5f465e076e902;
mem[751] = 144'hf727e37e0e80053114caf1b9168811680d1a;
mem[752] = 144'h1fbd165001181a59e6e11d961024e29518b9;
mem[753] = 144'h1c381b1907eceefd1ecef106e69cf193f858;
mem[754] = 144'h1ab2f4e407f0e9451956fbc206fb0a3f0341;
mem[755] = 144'he45a1ae0fc9bfde8f1f7fc0ee39006bdeb2d;
mem[756] = 144'h10c51a401bfdfedf192a166cf1fee771e450;
mem[757] = 144'h0ecef019f19be8e4e30b1a72e44de3f2f5a2;
mem[758] = 144'h1153e0d0eeb8eff4f81419fdeef6f0beff28;
mem[759] = 144'hf7da1da4e248144efc4e01481abe098314f0;
mem[760] = 144'hf696e0371188e0cf111be04e1c99f4b1fffb;
mem[761] = 144'hf0d406c6100de3eaf9c6e670153e068b0037;
mem[762] = 144'he84b1081e3c40ecd0c7418bf046f0c58058c;
mem[763] = 144'heb48e3ac1404e9b8e07cfbeb1b8df9c21695;
mem[764] = 144'hf7fbf93df4efe56fff95f970fddbef0ce7b5;
mem[765] = 144'hea681406edf7f976ee0df66802a9f13ee5ad;
mem[766] = 144'h1b111167f8d50a320a97ed61e30a18bbf43b;
mem[767] = 144'h088b10d21e0def8cf73f1491f9d8f640eef4;
mem[768] = 144'heba0fed11ff519dd09b0f95fe6601a4819e6;
mem[769] = 144'he2ed0bf01a9afcc50d3f175303410e4cea98;
mem[770] = 144'hfe1de8c7f2edefac06e9e696173e0c2b1ad6;
mem[771] = 144'hebd80dd0e9c7158deb841a2917b9efd6f6bf;
mem[772] = 144'h10a8033eea36e3ce084801a317d215daff66;
mem[773] = 144'he7930272eea71db8e07607eaf29006cf02b0;
mem[774] = 144'h03a8e0b213390207e209044c0a60e733f00c;
mem[775] = 144'hf9d3e0e3001c006309daf77bf597e1f30dff;
mem[776] = 144'hea21faf80809f1fee2f8121aff2405ed10be;
mem[777] = 144'hf4eefba6e95702371c2ff07303550e24e48b;
mem[778] = 144'hea501ea8ff80165f078504a90238eedcfae5;
mem[779] = 144'hf94f0c10f7d1e5f4ee79fb03f3a819ed1767;
mem[780] = 144'h1bbaf17b1173efd60e71f839000ee2d4027c;
mem[781] = 144'h0ac8fd87eb95026917e6e027ec6ce2bcf70a;
mem[782] = 144'hf60e0bb017920a6a0c311fa2f0d01321e763;
mem[783] = 144'hf6bef253013814591212e5c0fca1118c0a4b;
mem[784] = 144'hec8af711eacdfe3a1f0f16a0e46ffdccf7bb;
mem[785] = 144'he76008bf1a10ef4606bcf037e065157ceffa;
mem[786] = 144'hf13ff8a0e4c8f841e0ecef1df85d16a3e5c3;
mem[787] = 144'h1132ff4618b8ee1fe826155a1e3af29304c7;
mem[788] = 144'hfd67fb7811e7fd761b251505161ff86c064c;
mem[789] = 144'h1e56ff3701290e1cee14fe08ec9fefccf00c;
mem[790] = 144'he605fa771035e4b60e0cfa210914ffabe9bc;
mem[791] = 144'h03c1e2631b660033e7941b1cf4f91fa9e2b0;
mem[792] = 144'hf7af10f7137ae4d8e0cbe0caeb8919870aa9;
mem[793] = 144'h1e98fbd9f8f8ff2ee0ffedd1f7450f050625;
mem[794] = 144'he08f1a74ea8dffeefa2e06e7f0fbf2970269;
mem[795] = 144'hfa97efdc15d3f92cef98110ce208e9aae34a;
mem[796] = 144'h101ce76ff3a9ecdaebc5ea77114a1d040d20;
mem[797] = 144'hf58ce620fbf0f8a7e8be1fdbf0f1e0d3e79e;
mem[798] = 144'hf624e909f67714ef1e52f2530a090f86013c;
mem[799] = 144'he8fd003de5ef1785ecfbf102e96c0528e248;
mem[800] = 144'h1e510299e9b1e7f4f79e03f8fdd2e5f9f549;
mem[801] = 144'hf3df0e050d3a1fa605591bfcf38ee99d19cc;
mem[802] = 144'h10d50402f2ccf14df6051e320feffdf2f07e;
mem[803] = 144'h1974e4ffe2021394e101f90ce77de13dfd70;
mem[804] = 144'hf895f98aeb5cf4661fbbe6d70978fd0ff75c;
mem[805] = 144'he7f7f37bf0631a7c0b1614bfea13e01ef78f;
mem[806] = 144'h0e9ff4ad1e6615f5efcce65b1661fe280796;
mem[807] = 144'h12de1d17efde0d310d920cd104e7049210de;
mem[808] = 144'h0f2df53e02cf0ac014c20b99eb6e10100797;
mem[809] = 144'hecc4e614fd621321074cf4e00b54189808ab;
mem[810] = 144'h0a6ff4cc129c0ad8f71901990127ed29f81c;
mem[811] = 144'hedb8e8041a3be4511cfd1d6c030ef5511d2c;
mem[812] = 144'hf59eff20ec28f1fb18b8004117090ed8f78a;
mem[813] = 144'h15f8e897e5a7f07ce1091c461da0e0f80118;
mem[814] = 144'hf33d0ebb0e88060306e117f3faa603b1f91f;
mem[815] = 144'h12d9ecd6f9301dbde262e9e20c1a08d91a6d;
mem[816] = 144'h07cbfa1ee172e5081e62e77e1a791eda0b0a;
mem[817] = 144'hec2ef7a7fcd412e4047717ce1d9ce0e9fca2;
mem[818] = 144'h116b0891ef06edcc02280cbbea07fd58fb55;
mem[819] = 144'h012b01ede76defe910330efa0088f63a155c;
mem[820] = 144'he6e0e40d138a1a40e99b077f0e51e4bb0c11;
mem[821] = 144'h19b6e905e1090e96e870f736f2f411091662;
mem[822] = 144'hfae3f60ee71c1016fa0802cf17ee025016f4;
mem[823] = 144'hf10bf7e71af40255e6971f680c0b142eebb7;
mem[824] = 144'he1ebe09deff30832156c197f06410e17ec22;
mem[825] = 144'h135ce3cdecbd0b57ea29f68a11011642f5cc;
mem[826] = 144'he964032bf015fb87e0d40927176d15f6e794;
mem[827] = 144'h02cbe67205dc112fe2e40d3b0156fc11f77a;
mem[828] = 144'h122413781b421d170b8ce94de69efd71e62e;
mem[829] = 144'h0e38eda311020b7f0c90054af04be664063d;
mem[830] = 144'h0c700364e0a0034beca0f7a6f12f01880a0b;
mem[831] = 144'he9841469e1430e61f6861f4a1d1e15ae13b5;
mem[832] = 144'he71be4bd0471fe4de8d5026e007d0389e52d;
mem[833] = 144'he5e30846fef61614feaaee0efcf814b5f787;
mem[834] = 144'he15d02aaf623088f082d0a34e3b8139704f9;
mem[835] = 144'h160e0aa1f00e1fe40051f29a105be9131430;
mem[836] = 144'hfd260dd603fe1977e1960447f112e19c16d8;
mem[837] = 144'he512f5e51e7fffdd0d140aacf07bfb3a1761;
mem[838] = 144'h0aefefa10ddceb8214d4fc2c1c991bc91906;
mem[839] = 144'hf73e0564e9b91a06044d1e040812f4360627;
mem[840] = 144'h03e5188c194ae5faeb2b1d8f1e62e88ffb1e;
mem[841] = 144'hfd4717e2f4b70ca8f8651613fd96f19dee9a;
mem[842] = 144'hecd61674ebdcee6f1dc6f2a21e2ce6191e11;
mem[843] = 144'hf6ee048d0723ee5a147410b5125be1901ff4;
mem[844] = 144'hed7d1df90466f78fe7b1f66801fb02da087e;
mem[845] = 144'h1e14efd5fc510e32026df7ffe3f008bb0566;
mem[846] = 144'h1087012dfdb5f8511a9df8f7009bf69209d8;
mem[847] = 144'hf1d91fa9f5e20da91d9807c1146d041f19b8;
mem[848] = 144'h02750e171307e11c1092159f1d60ff57fae3;
mem[849] = 144'he36e0abaf5db121af073e301fba602ce1204;
mem[850] = 144'h1852f429164e132ffc97f4dff5be14c91992;
mem[851] = 144'heea406e5109e1c070e37f2b2e70afa57f4bc;
mem[852] = 144'he96c0e13fe1609ad1a52f0b3e7cf1d8319a4;
mem[853] = 144'h17f115b3198608caf8a2f64aedd91f55e4be;
mem[854] = 144'h13a1fa2f0a9014be0420085b13bfe3f4ea00;
mem[855] = 144'he7b704dceeb61cbe0f30e5ef1b81e736065f;
mem[856] = 144'hedf7196b16b00ac81270eefc1b5d11a51d17;
mem[857] = 144'h04a3eaa51d54f6c6fb2fe6f3077bff8af76a;
mem[858] = 144'hf17b0e52f3a6f318e8fcf4ce1794ec351070;
mem[859] = 144'he4480d7f06d31a3e137312430aa0ed2d02cf;
mem[860] = 144'h11c6f933ed3bee4c0a75e0321fb90e3900b3;
mem[861] = 144'h039fefabe825f1b8ed05f910f4f1e30def73;
mem[862] = 144'he73411c71b97e4bd077dee33f167f79f0701;
mem[863] = 144'hf26c14970a77fae0ee5ffca11db415e0e171;
mem[864] = 144'hf934f91ce3180a1d107e0324f55ee8df15b4;
mem[865] = 144'hfc84e66305f7f2c3fb041a160b511b5502eb;
mem[866] = 144'h1315ea32ea43ed5813e9e145144dec30edf8;
mem[867] = 144'hfb6afada197e037410b6f2ffe22be9ccfd93;
mem[868] = 144'hf2ca0f6ff704efbfe979e026e9a8ea231ce5;
mem[869] = 144'h06b608591de2ff04f737e85c01abe47f1c80;
mem[870] = 144'h18f2e399ec4de2390574ee5ae4e9e61e06db;
mem[871] = 144'h0127fabf15cf069f1af0f7bbf569e3dd1630;
mem[872] = 144'h1ac4e55405f4e74cf3baf8850378064ee8be;
mem[873] = 144'hebe9e92eea85038c0bbae94fec95f7c8e26c;
mem[874] = 144'heddf0ee918061facee121329e36010d6040b;
mem[875] = 144'he293041f1a29ee22f399e7821f201ebc139c;
mem[876] = 144'h1062e865ecd8125813e5f0540d59e1d4eb8f;
mem[877] = 144'hfa1eff38f225e189e21803f80dcd1ab5090e;
mem[878] = 144'h12a1f0391070e43eead5f154126cf9fff48b;
mem[879] = 144'h100805821d0e15b4eb1ce7960124031c1956;
mem[880] = 144'h0d490806f1691022fd01fc73fbd2feb0e545;
mem[881] = 144'hfb88ee07eeab1df800e416e0f02be526fa68;
mem[882] = 144'hf4bfe9c4ea1a195ce9450483f82ae1a51de4;
mem[883] = 144'hf792e717ee4d1a6af137e196fc3b150f0b23;
mem[884] = 144'hf8590c1ff7cbeefae5c2f2620abf1bc1199a;
mem[885] = 144'h163eefbf15e7fa331d8cfdcaf489e7f8e0ec;
mem[886] = 144'h0ac41c84f64de0b6f2f708a1f333130c14ec;
mem[887] = 144'h12e501e4120a0e6d184301edfaad182f16ec;
mem[888] = 144'h01270fd5e34c086d1b7f04f4f27b1f4903b8;
mem[889] = 144'he7a409ee0db501e5f8aded260b4c10f4eb6e;
mem[890] = 144'h05a61c40e5f2147af415120beeefedc01ad8;
mem[891] = 144'hf04ee5be15710220f69d16c30c41e725123e;
mem[892] = 144'hf4b0115df43bf9d50507fd970dc4e0e01124;
mem[893] = 144'hf8b9e23904880b7b199c1ea9e328f917e09f;
mem[894] = 144'hf15e065212060f6df68b16bde9ab14f6f902;
mem[895] = 144'he7941948ea8ee09d0af2fd1af2a902cd175b;
mem[896] = 144'hf540ff11f67de889f2c41b3af00418ceed76;
mem[897] = 144'he08fea5c1ca71f200ff903dcf52af6e5fcd9;
mem[898] = 144'h0ad1e8c4008e0fba1e63e2531e3fe3a3fbc6;
mem[899] = 144'h0c8c14430b1708abec601abce84e0f4e0618;
mem[900] = 144'h1b2cf0aaf881031a0dce1490f58aef27e06b;
mem[901] = 144'h0dc5fea0f861f183e597e28ef2381dfae510;
mem[902] = 144'h150ce257f8d90d89f2531dfae6ba007d13a0;
mem[903] = 144'h19d0f7b90ccbfb58f7b2e528f57ee4e6e9cd;
mem[904] = 144'hea09e129ffbeeaf41856143fee6ce0f5e2f9;
mem[905] = 144'hf0afe57cef07f893f03ee2f1ec94137ce78b;
mem[906] = 144'he9150b1608bff40c18f508521eebe2ffe9dd;
mem[907] = 144'h0e4fef71153cf5f3fb6c0c60033002c30a94;
mem[908] = 144'h0273e7a8189ef26d046b08a20b810f79f483;
mem[909] = 144'hec9f0e3f1d85fb641c2508810284f2d918da;
mem[910] = 144'h012ee9c3052c1199076ee130fc0013acf160;
mem[911] = 144'h1ea50e09f54601d4e0cd0a240e0a1ae6f7e1;
mem[912] = 144'he965f6680b21e8b707141f3a1eb50fc51749;
mem[913] = 144'h136aecdeeca6ed02f109f973e134ed3f0fd2;
mem[914] = 144'hf2f60d6d069c0254155cf0f106bde925123a;
mem[915] = 144'h1c71eff4145511d1e4100bdd1e2fe652e86e;
mem[916] = 144'hec61e0a1f067f924eb33194a0788e4d5e2af;
mem[917] = 144'h1d6f1f8ee5841808f07802c1e4e518240ffc;
mem[918] = 144'h1df001b4047c19b4f13c0c260cf9f836111b;
mem[919] = 144'he8fc15ae162be07c0d390d0bef3100350f0f;
mem[920] = 144'h1519e5131017f361ed0e182110f714e2ec37;
mem[921] = 144'h078c11ab13c40f9e1140046f0433056a0c0f;
mem[922] = 144'hf3b1ff40ea321beae73dfcbdfc6ceb6cf5cf;
mem[923] = 144'h1610088afd6affc014c21f6d0830037ae611;
mem[924] = 144'hfe7207ac0e0cfadaf092fb93069ff555e604;
mem[925] = 144'hfc1417090b15f5c61eb512290561ff1302f2;
mem[926] = 144'hf23903de1e9becd1e5fb0da40746079be581;
mem[927] = 144'hfdf40a4fe15e1654102c1adb1b24e3e4fe48;
mem[928] = 144'h1685000f19511178f3a9fcef047f124f14c8;
mem[929] = 144'hf02116bce1320bcce5a4feaa1b250933e129;
mem[930] = 144'h1b84fdc0ea541e14f5c4ec34f5a6eaf8019d;
mem[931] = 144'hedf200961cba044cfb2aeefc1c2b1485e13e;
mem[932] = 144'h09ecf6681e36104fea391fbb119f0b0b17bd;
mem[933] = 144'hec640e820eea19e2fa891da118a5ef5ef7d1;
mem[934] = 144'h0ff4017ded1503080d1818defcf8e7371817;
mem[935] = 144'hee830534e82901d1f873f639f999eb131772;
mem[936] = 144'h1016f1f7196bf56502baea75edd1e91700c0;
mem[937] = 144'hffd2018112320b7debc1165f1cd60b790e5f;
mem[938] = 144'hffb9f5f5e5980cefea3ee0c1f24cfbfafeaa;
mem[939] = 144'h11991cb7e885f1bc0a3118561e0d0429e82d;
mem[940] = 144'hff36067c01a7095b18521a84fc27e9b419b7;
mem[941] = 144'hf26bebe1009be628e6ad1c1be715fbfbfa7f;
mem[942] = 144'he8bd037a171ae27316b7eb57107d1f53e4a9;
mem[943] = 144'hf68beab914af0664ebace4a9ffeae8980e20;
mem[944] = 144'h05b5f80ff6dbe35e07fffacf1e111ac104be;
mem[945] = 144'he474039f0143fc1f081a071af882062101fc;
mem[946] = 144'hf20ce74008ab04270770fcc11b64080ef534;
mem[947] = 144'h1031137717eaec450ce7ffd11bb8ee89e801;
mem[948] = 144'hf93b195b0a47f920fea7e08a0ee8e566fc71;
mem[949] = 144'he4cfe1d10b55fd6f0cd0eba7e8ce0101ed60;
mem[950] = 144'h052be4d7ea6414f7eec31ac4f65f094ff952;
mem[951] = 144'hf3a0e793ea4dedbdfc7ce7301d09e5ae1caa;
mem[952] = 144'hf5d90b26e51d162d0e8c02e1fc671c56faf2;
mem[953] = 144'h1f34ef560f4e05cd1fb1f42e1d8aee4fdff4;
mem[954] = 144'he08d179210c2172be35ce7d404ef0ce6f166;
mem[955] = 144'h13bb0cee0ba1e985ea3517ede7ef19d8fbdc;
mem[956] = 144'he67deee9e403eae70ff10eece94bef200d21;
mem[957] = 144'h11641df80eccee2b03c5e8a81c96e36e0caf;
mem[958] = 144'h07b8e8e6e2060877e783f74cfcf8eb950ab8;
mem[959] = 144'he550f90ef450084f101a0ee40843ef86e945;
mem[960] = 144'h13b506d81d4bf8bfe7f90615fac6ee61e358;
mem[961] = 144'h1b72fbfcf34cefe5fc970a80fbce193ff9aa;
mem[962] = 144'heacf0cdb1603edeff37111321980e1e4fb9f;
mem[963] = 144'h014500a1f9321a001e8c12981ef6e6d8ee4a;
mem[964] = 144'hec620f910057f0fd1cb80ee70f1fe3fbfc53;
mem[965] = 144'he562035ffbd9fad80fdfe2af0aa4e50a1585;
mem[966] = 144'h1cf5eecd1aabf6c903cb1c75138bf0ae1590;
mem[967] = 144'h003c0df3ece8ebbbeed91c48ec5ee54af887;
mem[968] = 144'h07c4f4780075ee1d133ae1fbf67af5ed1b6e;
mem[969] = 144'he928e8350f85e497f48fe12911f9ed910a9d;
mem[970] = 144'h02c2f5e20229e714139e107019c6fbf217df;
mem[971] = 144'h1c9ff9e3e56df288154a1d46f470f7571219;
mem[972] = 144'hf2e5f41fe37e17e2f00c1ae0f6ab05dbf702;
mem[973] = 144'hf939f53c058fe69afc1509e70d13190efda8;
mem[974] = 144'hfdfc06baf2870549013b15b5ff8c04b90baf;
mem[975] = 144'he0a0028f0173f6600c310df7030b1a7ffa49;
mem[976] = 144'hf7c1e90c1fe7ef391f9af5b9ebca05caf88d;
mem[977] = 144'h11b0fc7218d7fb78004af94ef957fb19efa9;
mem[978] = 144'h0fb1eb85121116e6e5b608301672fe3b0df2;
mem[979] = 144'h10a5f3601bf700f3034df8560c5b0a6bfcbf;
mem[980] = 144'he208f2d1ecacf6330f6ee56ae3d50c7ef529;
mem[981] = 144'h1d8208e1e92a0349e265fc87e01508ae16e7;
mem[982] = 144'hedc0f8baf6bbf389f4e5015ae3aa01780807;
mem[983] = 144'hee1ee59a020f1d07055fed4506edf04ae5fa;
mem[984] = 144'h0721e2a8e116142a1666061dfaf306ba06df;
mem[985] = 144'hf6a8e7c7e587e999e7b9fae4115f0be71cc8;
mem[986] = 144'hf90af66f0d52eec9147efc41f9d5f54bfb70;
mem[987] = 144'hef6be9bbe3dce46f17e2f636f7381b4cf122;
mem[988] = 144'he99f1a1afc1c0db4e9c607f8ed84133bfe10;
mem[989] = 144'h1fb5e189e0dd019e027c0ff6fc8b1f7afcb1;
mem[990] = 144'h02150e77e2de1cc5ecaa15b7fc130e8419e3;
mem[991] = 144'h003c0afafe79ef87ef0204c40d87fdcb0f39;
mem[992] = 144'h09440664ff581d69f788fc04f10b1986e2cc;
mem[993] = 144'hfd37e8c10e4a0f75116f04c7e004f28eea30;
mem[994] = 144'hfe89136ff0ef172b0160f424f06f0b6b1aa3;
mem[995] = 144'h18601729fbf61fdfe2b7edfd0cf51d17023a;
mem[996] = 144'h1351ebcce6ae1bcb0b080889ee88e0211c23;
mem[997] = 144'h1dc6f834f3b7123e11a1f95a18f6076a1155;
mem[998] = 144'hed26fb53e428098af114ebbaec0ae24bece3;
mem[999] = 144'hf7e7f124181c0fa0e0e7e097e9e305ccec6a;
mem[1000] = 144'h06f90ac4ec7f043ffdfd18ef1394e43cf7fe;
mem[1001] = 144'h01d9e2e7f378f434117b0bfdffe718d60a4c;
mem[1002] = 144'h034cee50e7b9fe69f6440d88fd2dff191010;
mem[1003] = 144'he541e9bb0bfa03cbe80af6090dd8fa91f4db;
mem[1004] = 144'h008701ac0353ea3c02d0e659ed310735ec89;
mem[1005] = 144'hff0e024af90fdfbd108111a509f6e8d517b6;
mem[1006] = 144'hfc6d1cc007f413b1e70f1f9ffeb3e3ecede5;
mem[1007] = 144'hfce611221184173b0564e3670bccffcafdba;
mem[1008] = 144'hfff3124b0188f97c061de48a1cadf360f9e2;
mem[1009] = 144'h0ad4e9c61fa0e467197e08ac061001f7fd91;
mem[1010] = 144'h09d200e5f424f40d14d2f2b1f246e75918f6;
mem[1011] = 144'hef33e3acea67f82605420e40f7c414221f62;
mem[1012] = 144'hf40eea6e18dcf7ede4811387fdd8ea0a0d9f;
mem[1013] = 144'h1babf0530b89e3c2f4491e17ffe50b7cf647;
mem[1014] = 144'h1f10115aec7ee398f0f61472f1e41d65f7f8;
mem[1015] = 144'hf871e663059fefb5fa261797f06ef1d1f719;
mem[1016] = 144'h062504adf7f4059d1752fec7e1f512e3e3c3;
mem[1017] = 144'h0bd81295fd4e17e21d96e966e727f033e191;
mem[1018] = 144'h09aae458f8431ac11fd11d54e092e0b418ef;
mem[1019] = 144'hee1809f5017a02d0e69e189e1313106d1ae3;
mem[1020] = 144'h073413b3e1f5e59815270fbc0cb0f8fa1795;
mem[1021] = 144'hfe3cf50d00c9ed7cf99ce57cf8bb0ceb1e8b;
mem[1022] = 144'h13b714210a270881f8a309ebfb3a1974f6b7;
mem[1023] = 144'h1c9cf20bfd10ee33f0ca0fece8ebe26e0aad;
mem[1024] = 144'h1f7d0ecb0c8311e41dc2eb80e44cf80bf165;
mem[1025] = 144'hf391116f0a6019acf1b9fb6dea1bfea10f40;
mem[1026] = 144'h1ddc031aebbaf4ed10e4e50211ebef1ce89f;
mem[1027] = 144'h1c240ec5f3d8ed38f1d8117ae41a07e40dec;
mem[1028] = 144'h0fcee4daf73bfee2f397151e1989f1931c17;
mem[1029] = 144'h0bf603bd003dfe34fa8e0ae11bfe15bd1df4;
mem[1030] = 144'h0110169d0064f5b6004fe32510341bb00d9e;
mem[1031] = 144'h0f1df96ef4dbe6cbf88d0b6f132deef11b3f;
mem[1032] = 144'he1e5eb740e990abc08a9f0cceef0f1cd02fa;
mem[1033] = 144'h0105e50502db12cdf92aefa91a99162be34d;
mem[1034] = 144'he48d1c0205840676f1cef05b1edfe374eefd;
mem[1035] = 144'h1e8ae2511ae1e1420c4e003eefc41f4ffef6;
mem[1036] = 144'hfbb7055d0b19e7a4eec2e5e5eb8a051e1998;
mem[1037] = 144'hee18f03de26cf64cf3bcf514ea9c0be70665;
mem[1038] = 144'h0a46fb8002ee1f651d91f311f194f4e9eb23;
mem[1039] = 144'he42f1f9c08930cc1fd4c01910e4c18800186;
mem[1040] = 144'h0df5f72f0ab4fc62e3fd1e2a1ece059bff93;
mem[1041] = 144'h06901ea10ad3f7a4e402ebb81e5fefb01b29;
mem[1042] = 144'hf408ed4dfca315c31ca6eb010ce4f280e7ac;
mem[1043] = 144'he1bd19a80b950eb002ad0c5cfc61f5011eb7;
mem[1044] = 144'h05cdfbf7fd09ef3f1bf5044d02d5f42c01fb;
mem[1045] = 144'he8da104d0f1d1148e5cb0eb3e1161129f4a9;
mem[1046] = 144'hef3c1c86f95d17fe0443e862fa050151e17d;
mem[1047] = 144'h13df09c60bf51ffce930eafceef3ed26fc17;
mem[1048] = 144'hf8c701de0917ea97ee35eba71a17e20e0194;
mem[1049] = 144'he5cefd8ffb430ae80b52ece116bae7fffae4;
mem[1050] = 144'h13e8f33307c1f044fefce718198bf6dc1362;
mem[1051] = 144'h1a53f8f6fcfe171be3951451f044fb89ed47;
mem[1052] = 144'h1537f5ab0f471fc2e5dcfbdcfe36e2ef1df4;
mem[1053] = 144'h0402e4a2ff15e23a03080299035e1b6a0756;
mem[1054] = 144'h1fc1f959e143fc8d0275e281f73303981816;
mem[1055] = 144'he2731e971453fd7f07bde39f070bfaa1e791;
mem[1056] = 144'h096618a106961d83046b03691d851c131e83;
mem[1057] = 144'h0ac9fb70eab602031b3612450a101ce81a5b;
mem[1058] = 144'he4e41237f4e8ff86f5590e29ff85eb0e192e;
mem[1059] = 144'h03f0fdb31bc9f410fc5707a902c0f1c0e374;
mem[1060] = 144'hf2f9f162e426020016d8f0a5e3a80db3e165;
mem[1061] = 144'h0975e62c09820d47f653e7080ca0e37d0418;
mem[1062] = 144'hf8b5e79319edfa67e7961baff4600825f22a;
mem[1063] = 144'h10131c65e4d80a760f5eeb4ef7adf448f82f;
mem[1064] = 144'h1c691ccd1ecbfd23e8f3178d15c814601954;
mem[1065] = 144'h1d5f169dee67f9c3f2faf0ffec7808d0e934;
mem[1066] = 144'he4991afbf0c2fc5e1220f8f4fcfb11371d88;
mem[1067] = 144'h086d0bdb1252fa55f85a16021e3e06391840;
mem[1068] = 144'hef47e38b1c48074dee7a1ed7156401cb1286;
mem[1069] = 144'hfeafe5981ba31d20fa8c04961874f22e0c05;
mem[1070] = 144'hfb3df5cdf0a51cc10bb303ea04d11b19f44d;
mem[1071] = 144'hf1d81893fb73eec7067b0b5c0b77eef918cb;
mem[1072] = 144'h152e08dcf8f1fd781df4fda7e0e1e02405c1;
mem[1073] = 144'h1d4300200c6e18a8160f01a602b1ed58e18b;
mem[1074] = 144'h12a701b2f1e9e352f8f1e5ba1deef4b809cc;
mem[1075] = 144'h18fdfe0a1ca2e786e78010ca0292fbcd08c3;
mem[1076] = 144'h1431ef2d1673ed731904123612d904981481;
mem[1077] = 144'hfa14fab3e4570b49e848ffae11d0e53fee2b;
mem[1078] = 144'hed9fec04ef8f0022e320f1fafc12161e07d3;
mem[1079] = 144'hecf7effdf261fe0df4c91956f4511c37fe62;
mem[1080] = 144'h0a391ce3f8ddf708e9461aa5153811940f0a;
mem[1081] = 144'hfc9009d2f6cf1d0aeeac087af8431cb5f548;
mem[1082] = 144'he6c4ee2e102fea80ea49eff6e0220751ea70;
mem[1083] = 144'h1f821cfef844ee9ff1c706c11e20e86a0807;
mem[1084] = 144'heca6e8f908d1f11d1f5c192416b8e04d1338;
mem[1085] = 144'h0b8900e5ee5e0beb01d81831f8a7fce8e01a;
mem[1086] = 144'hf3f50481edabfe971b4e0b970be7f837fbcd;
mem[1087] = 144'h017818530fe915adf3a4e33201cdfe141caf;
mem[1088] = 144'hf81cfc05f88af19f0df5f8b51ce81864e4ca;
mem[1089] = 144'h18681fe0edd403b705241ddef63601eb1807;
mem[1090] = 144'he8dbf61bfd85f956f4f006b70eb2e58e079b;
mem[1091] = 144'h184def930e6015d01678082f00d31af8e692;
mem[1092] = 144'h036d1c6b015f0708ef5c000ef439f0ece37e;
mem[1093] = 144'h0db91f2e2172f7f10010e0a9e531200512a2;
mem[1094] = 144'h0338f842f2060486122010d7039800bc191e;
mem[1095] = 144'hf52f16610c6618a714d1fb36116ef4c9009c;
mem[1096] = 144'h1b831e251548fac5eae7fb50fdc1053fe52e;
mem[1097] = 144'hf8c1146d1afee4e0114df01a0fd20e0f17ec;
mem[1098] = 144'he7f6e726f83c08911a17e4bf03c4ec5407b6;
mem[1099] = 144'hff38eefd0fa3e6170faefaa41a85f8ad02d5;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule