`timescale 1ns/1ns

module wt_mem6 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'he735f53e0fdeffc80582f0ac1de2ef040143;
mem[1] = 144'he5671326eba3f994fb90f0e2f0a51a4ae950;
mem[2] = 144'h1454f83bf67212de13f01c15093c0219180f;
mem[3] = 144'he6d511dc190509d70dc3f563ffa119d70cb8;
mem[4] = 144'he352fb0ffabb0f3903111eedf13a1c58f34d;
mem[5] = 144'h0dfaf4cf11d81dfee6c3fb1a0201071ae5d0;
mem[6] = 144'hef1ffccf114ce7a4fd5af66606de0a550a45;
mem[7] = 144'hf14cfb841139ec9c18d1f9651497f90913bf;
mem[8] = 144'h1135051e1735052ee114fefe1b67e7ba1610;
mem[9] = 144'hf644eb561981fc8c0a6be790e379f52c1f42;
mem[10] = 144'h069f0d440c5201ac120203a00eb4f26ef961;
mem[11] = 144'h0c7709f4ebff1085e706f109fbb01bc31310;
mem[12] = 144'h01f6f576fb0d1546f326f704063dfcf703bb;
mem[13] = 144'hf451168b1cdb1421005cfc6a128008afe3d7;
mem[14] = 144'hebbc07a7fa55e2ab1c211effe6d8f6af1c84;
mem[15] = 144'h00a6e68000151a02f904fba10840e37f1fd8;
mem[16] = 144'he29b0a49f6ac1e44054e0773ec170b2e13ef;
mem[17] = 144'h063e0325e1a818940e9efc941c6604ea095d;
mem[18] = 144'he782efbf02fc1423f5ec03f4f4c9f809f952;
mem[19] = 144'hf8bbfb8a123111a30c660d280efe1c7ee6ff;
mem[20] = 144'hf336f9d5e8faf9b0f8f9f0a51556f712e58e;
mem[21] = 144'hf9d90360ef90031cf196e9dee31fef751d36;
mem[22] = 144'he8640756128bfbd8e0b4ef10e5db04b2fcab;
mem[23] = 144'h14e7f45c048b0b52e890eadded490af9e973;
mem[24] = 144'he34b01f9fba3f37a19ad02ba052102980d97;
mem[25] = 144'hff4a025bfd85ee1a10c608ebee7af63f1ab6;
mem[26] = 144'hfa01e9e8f03ae257e93af4c10fb906c9f9b8;
mem[27] = 144'h1202191bee67f782ef87f6670face84bf260;
mem[28] = 144'h1da8015d1893e57fe5c4fc14000819e61207;
mem[29] = 144'h1061e74be33e069c1ea1fdd61221164ff4d7;
mem[30] = 144'hf6261d0f118f1c91e4b61a4b0135ed36120f;
mem[31] = 144'he3750650078be152e74ce47e0b9d12f6e46f;
mem[32] = 144'hf3fdf9f2e6c90c68f2e40601e5e1f39ef217;
mem[33] = 144'hea09193ffa2bf4deefcf0d50f41af3e2e931;
mem[34] = 144'h0182f86c15f3f31f045419850d0c18cd1c14;
mem[35] = 144'h1d4f18b81428e61cefcee8fee247e0921850;
mem[36] = 144'hf5b7f9830aa7f2590c7cfc52eaf0ed07fbb5;
mem[37] = 144'h17ff1996fe5ae7bfedf2157116cee4edfe0b;
mem[38] = 144'hfdeb0db009b8e90cf3b401f7e45c0af40dc4;
mem[39] = 144'h059f0bbbfa00e92306f30850e358ee0f038a;
mem[40] = 144'h0829f8ef06731a750f61e5730a7c14561b0b;
mem[41] = 144'h0f03e7b6e16f08ca1ed3e372e4baffcce904;
mem[42] = 144'hf1c2fbf7ef85e064f37a1bf3f7fbf29e170e;
mem[43] = 144'hf6781f8c1a6de37aea66fed30d5be7451684;
mem[44] = 144'he719f5e50151f80314551196f524020de7b3;
mem[45] = 144'h102fe45b0302ffca1dfdf9ca175ee652e6da;
mem[46] = 144'hf6961ce8f708f62ff30b0f67f038ea1b0d25;
mem[47] = 144'heeff0761f234fdbee7d90f1607a4e7ecfa53;
mem[48] = 144'h13ccf117ee8706ecf076e319fe9dfeb7ead0;
mem[49] = 144'h1cd6e56ae4aefd7b05420528f269e9ccf25e;
mem[50] = 144'hfd5feaebee730560f991f717f5c71ae0f4b4;
mem[51] = 144'h048500e0ff9c0406031a023feb4eea94ecb9;
mem[52] = 144'h03061f111a1b03690896047c08530668f573;
mem[53] = 144'h0eadeb8f19fd170804b1e4f30820ea78f5ab;
mem[54] = 144'he764150e09e5e525edbfe1aef711128f124c;
mem[55] = 144'h1adaf12ae6ac091710e3fe11e6be138eee05;
mem[56] = 144'h1dc60792f25b0835f8830d32e8731f6f0241;
mem[57] = 144'hfec5ffd3f0cce442115d09ab1975e3dde88d;
mem[58] = 144'he172022ee9ade42af779e98d1b21f749f670;
mem[59] = 144'hf3f5e026efb0194a08f9e41b156d1367f0d7;
mem[60] = 144'h02e511c3f3a40c14f988e3ebe96f197cee0c;
mem[61] = 144'h12b3ed0beaaff5581d5cfc560c550d8f0883;
mem[62] = 144'hffea06be09eb0f4604e51835e0d913ad19c1;
mem[63] = 144'he4e41322099afa4b1b890b6de927e04df03b;
mem[64] = 144'h1c601b7cf0a6fb531b33125ce21ff6ef00c0;
mem[65] = 144'hffb70a1c07d4e9c004070dd1eec5f2adf1f8;
mem[66] = 144'h0dfbe45400750ad9e60104b2e56f068318c8;
mem[67] = 144'h0e2ffb36f397fda615810a901b0816611eaa;
mem[68] = 144'hf3bbe09c02cc13180f6cf2b00fc70c83fdb8;
mem[69] = 144'h1b8de817f14f1caa0eb0f57a1f7e081006c9;
mem[70] = 144'hefd8f0f3ee35f3c4fd7ae08bf9a40dda119e;
mem[71] = 144'h131beb620695f7fef41bea51e286158910f9;
mem[72] = 144'hffa7ec4519d2ec4311ed0631f255eeef1f8f;
mem[73] = 144'hfda3f32e0846e59e1833f2400c13efd510c9;
mem[74] = 144'h0c02fe06f77c1808fa8c1d9c1d96ee62fdf8;
mem[75] = 144'h057d0263f341edda03ac0743fecfe0e20bfc;
mem[76] = 144'he22de384e99417b0f99b1abcf1381ed2e64c;
mem[77] = 144'h1873e65d18d11617ebc1012513fcfb900e45;
mem[78] = 144'h11fa0f4f020504d5e2aaf8fdeda4e8610a23;
mem[79] = 144'hf35816f41d511a3707e819cafbd91d531460;
mem[80] = 144'hfa2ce6710b5a03a5ff79f022e18fe9d1e699;
mem[81] = 144'h1cad091c01c8f073e89215b5efa21a1def48;
mem[82] = 144'h1fb3f5c1ff17e3d51eb5fc1ced40e1870a9e;
mem[83] = 144'h12140a55f29c080f09dcfbc9f7e20f77f2df;
mem[84] = 144'hf5401031ea83008df11efbe8174b058a1842;
mem[85] = 144'hfabff8a3eff702960167eca6f890f252e3a5;
mem[86] = 144'he7301326f27befde1347f73aeb7f1965fc72;
mem[87] = 144'hed25e23bf7b11c0bf7901d8603a8e3b0f779;
mem[88] = 144'h15430067e6c6ef5bfd01f42afe55fd2306ce;
mem[89] = 144'hee7e0ebcef111f61e226fca8f74ae27e0a20;
mem[90] = 144'heab60cae1595fd5ae2e8f28de4a501b6001a;
mem[91] = 144'h1628e00aeb030879002f08950876082e1a7b;
mem[92] = 144'h123f0fefe5d00110f056e1e61f41f869e5cb;
mem[93] = 144'h0ac2fb981b4f001910aee4461cb7e5ad15ec;
mem[94] = 144'hf798e1a9f3bf06b9e616ee0e074aef1d16c0;
mem[95] = 144'h07511618e0d91f58fc13f5bdeefee7901039;
mem[96] = 144'hf25a17801c99f80ffa5fee851ad3e5b10b21;
mem[97] = 144'hf0ac0e41f5c6181ff140108114d11a6cf33c;
mem[98] = 144'he55beb551719f89809cde1c303c6f8d6e7bb;
mem[99] = 144'h1c4af4a2fb8d002a17a1e1f71f4f0a621ccb;
mem[100] = 144'h1b9f0d0a1a06e78cefa20b84e169187f0ee4;
mem[101] = 144'h14171dc21c7c0356095be4d7f5f8e887fb54;
mem[102] = 144'h0696f4641379e303e7260c231773e780e741;
mem[103] = 144'h09261851026c00bafd09fdb71e71f8caeb8d;
mem[104] = 144'h0f41ee5304f61140016f1856fcbb1c611bca;
mem[105] = 144'h1d180fcf0b0be5360fb71864095cf78ee447;
mem[106] = 144'hf293f8371f6e09b316871886ec6d0bcdf8a5;
mem[107] = 144'hef8dfb82e1dd101516a3f91b12baecadf56f;
mem[108] = 144'h08551bc600941e34160611f41c251f91ed2d;
mem[109] = 144'h1a881a70fde912e212f8e4d012a606f00d57;
mem[110] = 144'hf1f0fdc0fa0af5d3ea1407e0f5a808e80458;
mem[111] = 144'h1b9113c6fbb1159af5bde91012770001f938;
mem[112] = 144'he90efb3d06b20d53edf0fb96ec7f00a6f531;
mem[113] = 144'h0908f90e05d8e540e17bfd03f07f0327e60e;
mem[114] = 144'hfe01efc71e38ff58f23ee3500a59e3a00dcf;
mem[115] = 144'he314063f033712af1748fc5102c9e6e2eb19;
mem[116] = 144'hfdf4f6ce04a71813ea95f031165f1d4305b6;
mem[117] = 144'hfc2beeb8e9e1f27b0f831a980d48106ffe30;
mem[118] = 144'h1e070dc9187eecc4f896f9e618e7fbe61fb3;
mem[119] = 144'h0c741ee6f431f7f41afce54e0d5b01baffb1;
mem[120] = 144'h0078ffe1eface0101d111df71d3314861817;
mem[121] = 144'h06c01e3cf252134c0cc4131d05680a5fe777;
mem[122] = 144'h04400c34ecdd1fbb13cae919e01b0fa31a24;
mem[123] = 144'hf9d7e3f4f05fe9a7ee2cec05099413241889;
mem[124] = 144'h042ce403fc2009fc2087eb580114e517035a;
mem[125] = 144'h049617b8072fe9eee74dfbe918a9f3b9e467;
mem[126] = 144'he2f2e889fd0eec511905199e1fbae00b1438;
mem[127] = 144'h171be446ee7de773f1c20f1816a0ea62f56d;
mem[128] = 144'h1cc9e971112ff6e916b108f40a74189216e7;
mem[129] = 144'he477ef9a0984eeebe7a5ed04e7d51635027b;
mem[130] = 144'he6090e9710bf11aa17adef4d1c2a0c30fca7;
mem[131] = 144'h133fed80e7e10d7910c7fde604131588e027;
mem[132] = 144'he0010ae81619ed2606dc17d113b0170ce671;
mem[133] = 144'h10ddf2d2ef0c10fb17ea1d2f076f099bf271;
mem[134] = 144'h10131a91144ef31715f7ef2900b9160f0b6a;
mem[135] = 144'he66a057dec7905e30c0317341e141583094e;
mem[136] = 144'h1e26fbcf0e88e39dead51aec05e1fa97e5df;
mem[137] = 144'h14d7e4121b72ea4517f7e089e0840f2e1316;
mem[138] = 144'hf9aafadc0e9ae5d1013912481802148e099d;
mem[139] = 144'h0d5c082408cfe315f495eb3cec6af41d1811;
mem[140] = 144'h198ae90c167ef770fa5a0c2718d0fa5d1304;
mem[141] = 144'h1db21186f5160a6310f3e83df66efeb7f084;
mem[142] = 144'h08760ffa19df1b26ffcdfa34ff3de07cf48a;
mem[143] = 144'he1a70d84f3d4fe78e3ade4cfe54efdc004db;
mem[144] = 144'hfb06fac40a5b0ee21125180de992e2830394;
mem[145] = 144'hfd721a841d70002cf1eee0a40db3f1f8ff91;
mem[146] = 144'h0e69f272efcae976e1eee826e293014e0906;
mem[147] = 144'hfde0ec23e8590471ea94e0aaec07fd1d1839;
mem[148] = 144'h0e73e5d31e72f2af075d025102bdf481e166;
mem[149] = 144'he0900e720473e791177bf6ff16670108f15c;
mem[150] = 144'he72d0d070a261f55fbc01d3bee9d084dfc4c;
mem[151] = 144'h0f51f7a41700e4ef128fe1af19941b44f5ac;
mem[152] = 144'he394e06307e7143a0c04f68bff710dd5f21a;
mem[153] = 144'he99f15300d691d70ef6fe263e6aee52dfb19;
mem[154] = 144'he71ee06b1f18fa42edc8e40217101ae81649;
mem[155] = 144'h12e80cc5e62cebfa0aca140afd190669e638;
mem[156] = 144'h0235eb92e24a1903fe2eebdceddbeb250154;
mem[157] = 144'hf80de338080de470fd3e0b5819c5f5dce242;
mem[158] = 144'h0ee41087f132f334f3a6073715e91fea02d7;
mem[159] = 144'hf126f50d1386173012c8047cfd8d1e38f401;
mem[160] = 144'h19a1fbe4f236f0ff10b6e978ee4805e8169a;
mem[161] = 144'he806fbe111fc1cef10dc045214d3efcc0fca;
mem[162] = 144'h1a5fef300b47ff1310b30857ea79e4de0987;
mem[163] = 144'hf1dded55eea4ea0ee51605fdedca09a4166f;
mem[164] = 144'hf99114a612f8f29d1b5c1a65fbc30a78e565;
mem[165] = 144'h1faee92c0ac7ea94ee94e6031c5b0c92051e;
mem[166] = 144'heb3de58f1f2f1e4c1f6fefc71b5b147fe9c6;
mem[167] = 144'h1e761a54fcecfb190a9318f50521024f1fd3;
mem[168] = 144'he6ceec76fd20e8a6f6fae806ee3be1f4e376;
mem[169] = 144'h060c06f4fe68135014e002db1608eaadf788;
mem[170] = 144'h16571c841e4405131cdae002e14f16e70927;
mem[171] = 144'hf09315cc0f5ae349fafd11c1f374e26cfee6;
mem[172] = 144'h0bc316f0e5490dfc18bdef481afbfe9cf60f;
mem[173] = 144'h01421a59055409ade70ee5410be30a39e558;
mem[174] = 144'he2f4efd3f4731c440b2e1f3b12cb0f5c1cf3;
mem[175] = 144'h0e74fe3dfdee0057001006a3f1051e640bce;
mem[176] = 144'h11daecda0856eec0efcf1de0ecfdfafa196d;
mem[177] = 144'he3260c51136c0134e4f8035d1dc9123a143d;
mem[178] = 144'he587e8f0109fe4d71923fe84fc09f9ff0b73;
mem[179] = 144'he2dd0da8e6d7080b0090f34eff0e19e2f584;
mem[180] = 144'he178fb16037718071d54fdd2068e19f6fd21;
mem[181] = 144'he4c9160ef1b21e8af33d19131ef4fc5c0270;
mem[182] = 144'hf4b400710b170045f748e270ecdce4c0f3fd;
mem[183] = 144'h107108c703770fe4e38d13920d9efe311838;
mem[184] = 144'h0f82108711bff43fe51fef6c09631569e978;
mem[185] = 144'h1063f80ffa78e7c812f001abe9a416ee10e6;
mem[186] = 144'hfe901534e5841163e8f9f394e075018ee9aa;
mem[187] = 144'h082bf950efb5eac2028006c2e1e605b6e09a;
mem[188] = 144'h1d38f78a1f0601fd157ceb9819b5e51bf0b4;
mem[189] = 144'hec43f40be0ed0082e9150c791692e268131d;
mem[190] = 144'he5f51d9c0978ef310c3f0bddf15816791cdc;
mem[191] = 144'he6c2ed860d920d7619fce9b61a3ff8810875;
mem[192] = 144'h1b00e4610bd01f2105f1f62f11bf1a1ceb26;
mem[193] = 144'h189fe419e5090ddc08be1184060f0681e3eb;
mem[194] = 144'h0147ee2005841265079be70af4d8fb88e3c4;
mem[195] = 144'h1267f02ce5f41b41e5f414dcee0ce716e64b;
mem[196] = 144'h08d1e68017e1ea4e1351f7e1f5720bdeec0d;
mem[197] = 144'headb10f50186e449fa33f88719c4eb40f6f5;
mem[198] = 144'he58f11adecf205bb1158f0da0afc1eb4022b;
mem[199] = 144'hed38fe150c0d0389e41df8bc15ff00bd1c7c;
mem[200] = 144'he5eaf46af598ed18f2f2fedff5d11b6f0ffa;
mem[201] = 144'he7e314ff10f018081353eeefe74619911339;
mem[202] = 144'hf88b17a7e4adf4250933ef10f4dceb40e764;
mem[203] = 144'h0663e2870a61040c0aa0f3d5f43a1ed6fe2d;
mem[204] = 144'h0ed20392e24ee42a036b0242e7cee1a702d6;
mem[205] = 144'h0eedebefe122f528f97fef350a5d17fbe3c5;
mem[206] = 144'h07bdefdc1287f079e17ee75115a7f348e2f6;
mem[207] = 144'hf37ce96110c11ce10e8004fe16e30cbc05fb;
mem[208] = 144'h03dc1e8aec2a103dfe780772f6d0f874fb67;
mem[209] = 144'h0524171cfb75093af7fe08f908bfef591d63;
mem[210] = 144'h035a144f1483f92e0e15fbd2e5c00a2cee48;
mem[211] = 144'h1986f144ec0f1eebfc041a9e1bf106a20830;
mem[212] = 144'hfc1ee63ff1200e4207360c6211cc1ff2e4cf;
mem[213] = 144'h00e413b0ede4105cec35ea1ee2011cf802e8;
mem[214] = 144'h10f50028e93b0ed80aca13a7fe180e04fb98;
mem[215] = 144'heb2518901240e946ed010a040c041bfb1cb1;
mem[216] = 144'h086cf644e997eb4310161abd0bcfe243f969;
mem[217] = 144'h1f3af205f3641790e5eff7f5013f190bf9c8;
mem[218] = 144'hedeb1706fe07f4a6f9defdae135e02dff3f3;
mem[219] = 144'h17c20051f3f80adc009607531c5ce2effeca;
mem[220] = 144'hf55814a0ee721e400ec8f65509c603b8e5ff;
mem[221] = 144'hfb110993048dfc69e0930809092b057e088d;
mem[222] = 144'hfdf4189018aaf0021f87fcbffc7eea280e91;
mem[223] = 144'h101afb10e82bf8df0c411f4be9c1f2aeecec;
mem[224] = 144'h11d30f82f5a612560442ff1909e8e0781217;
mem[225] = 144'hee8f192df8be00ccf55a0e721dcbfac0e398;
mem[226] = 144'h0bd9f8351b51ef1dfdb019b813dcedfaeac0;
mem[227] = 144'h11a5fed50bbe0e48f3f7f11cf1c5e10cf9a0;
mem[228] = 144'h05e0e6cf1c3a138e18dc1071e631fff6f50f;
mem[229] = 144'h11dc19930433fbb0ec740915e58fe160e5d2;
mem[230] = 144'h00fae3bfece11fb6e8fa12fc15ec1ddb190c;
mem[231] = 144'h1a4beb7a132bec730126f5e3ea66e454e17b;
mem[232] = 144'hfec80b0207efebb9123af1c4199afc750cc5;
mem[233] = 144'he463e5f01c78fd3008830a4bfaa8f156f899;
mem[234] = 144'h04d2015c0ae5ebc1e198f1490205193cf573;
mem[235] = 144'h0ed7fe65eff7ee9c0ea1fcecef63e689e0dc;
mem[236] = 144'hf3e006151ac4e064134deace0014fac604ee;
mem[237] = 144'h005f1373ec76fa8ce43b069dfad7158c1019;
mem[238] = 144'hfc10fe46e24feab1ecbd13e0f9dc0311f0ac;
mem[239] = 144'h1cd210d80700eb0ae8d7e7631a5aec66fe6e;
mem[240] = 144'he391031b1e72eceefa8ef7d3e300fd92f3d0;
mem[241] = 144'h0de81dbc0fa3e6cf050203b60443e9e4128c;
mem[242] = 144'hf32e0a9808cee52810920437f992e5311b6d;
mem[243] = 144'h1599ee2002a8ec01f844f2f21d00e5d61b65;
mem[244] = 144'h078d07991f600f7a01351a24fcedf177ee8c;
mem[245] = 144'hf6f618b6f758e90ae978e275f71004a9f258;
mem[246] = 144'heab50ac0e6581ceee62fe81ee1a1f645e9c1;
mem[247] = 144'hf14113381bc31c82e5abedede8fcea65fd95;
mem[248] = 144'hfef5066bf1b41d4a0da60891f48013dbe59e;
mem[249] = 144'hecbc059aff62e2c41899e7f70c0a073def3f;
mem[250] = 144'hfe1d09f0e767e900030ae4181d60032e0e80;
mem[251] = 144'hfbc1076aee6f1dec16af06a504b008d5e778;
mem[252] = 144'hed2ee34612fc1f66f4cc06fe19cceef2ea2b;
mem[253] = 144'hfec40d7dfb55e60b1ff8f85108730bf80ed4;
mem[254] = 144'h17fff6eb0cf3e3e8ed6ce368f9b6fb731c3e;
mem[255] = 144'hf0041adbee23feecf2c4e319e350f061ef18;
mem[256] = 144'h0f841a43e8870f0ef4a70a56e2d20c771fcf;
mem[257] = 144'h1bce12251c03f61e1e2eed34e426eabff28b;
mem[258] = 144'h06851be4e132e50ee0750ebe09f1fdec00f6;
mem[259] = 144'hf60bf6b3015f170c1fb8e5eb142819f7185c;
mem[260] = 144'hfd10ecdd1ab612b2fda7e3fd10c40c61f594;
mem[261] = 144'hf2c6e0efff57e32a169fe43be7041faaff65;
mem[262] = 144'h0528fa3707e4e0461e55e836fce306440082;
mem[263] = 144'hec131a470cd0117105901648f61811720d52;
mem[264] = 144'hfb05fa56e10103cde64405cdf33ce49b0a68;
mem[265] = 144'heea10ff80b78e996f2cdff650d8c1434f521;
mem[266] = 144'h005be7b7e1bdeb3bf2811523e6eef431100c;
mem[267] = 144'h1690194b0230ea4419e6086d1a7af41c1e7d;
mem[268] = 144'h04e2105de64af8d218da033b130de3f8ebb0;
mem[269] = 144'h10cb17231518f54ff3691c44e67aed2fe46d;
mem[270] = 144'hf4f8e4800dd91650e99c07d5182fe99207f7;
mem[271] = 144'hf0d6f27c021d04ad0828e10d0a890a0cfd06;
mem[272] = 144'hf2a5eb7c135e0831f394f332e271e26ce756;
mem[273] = 144'hfb1bec1900200e9015ff1ab6e3450b42fe63;
mem[274] = 144'hecaafb3deba21b3cec6c1e9004470ea00ae5;
mem[275] = 144'hec3608cd1c44e83217a50e70f6580304079e;
mem[276] = 144'he324fb16e2620ca9efc21224080d1fae035b;
mem[277] = 144'he9b50323fbba1e241a7f01e8f990ea58030d;
mem[278] = 144'hed97dfec0bdd18a7e955e42dfacdfebc0e6c;
mem[279] = 144'hfbc512210e0a11950926e56b13ee0d69183a;
mem[280] = 144'h053a12d01e1d113afa5ffbd6e601f4f2f896;
mem[281] = 144'hf44cef9ff4011f26f04de57e1da40fc200c4;
mem[282] = 144'h00790d24eb7bef631b9418fe14890420fccb;
mem[283] = 144'hfa3b0dc4ff0b070cdfa60fb4ed20ec6106d7;
mem[284] = 144'h13580daaf30a14f81711ef35e9a2e054e9a7;
mem[285] = 144'h0390eb0b1540e63ef89ee001e9b0e29c1aab;
mem[286] = 144'h04eef6ace6dcf4711a581a72fdbcf45cfa18;
mem[287] = 144'h1243f434010af2671a0cf3e20322111e19b4;
mem[288] = 144'he193f94413a91cf105a5044a0595e4b10365;
mem[289] = 144'hfb89eb57186808cd1df91f00166b1966f6cc;
mem[290] = 144'h0a0806bbe1b6ed1ae5db05a2e033074b0ab7;
mem[291] = 144'hf8380ffc08cd0f951caa0debe162093b1936;
mem[292] = 144'h0e0f13c7058111d11083eabee018ed771df9;
mem[293] = 144'h19f011c71bcfeec211db1ab00f390045fad7;
mem[294] = 144'he9f20b25f478ef99f6bf151ee301152b0e8e;
mem[295] = 144'h1a6013f2ec750326f70219c0e04d0d9de829;
mem[296] = 144'h0ff70c10e75416221a75153ded03ed38fbcd;
mem[297] = 144'h0097f920f8a5ff7b03c3e03bfa0cede01bd6;
mem[298] = 144'hf4b4121d15bbf01e10a5e58a0c13ff850f5c;
mem[299] = 144'h13de1df3f2e1e32cfda4e2d3e8f5f235e492;
mem[300] = 144'h083e07540f381390005215d0e4a611d9e023;
mem[301] = 144'hf8b9e333fe65e3f2f3260e7ffa2afa54e2e1;
mem[302] = 144'hfa1a0604ef05e8cfebe9e2bf142e121ef3f6;
mem[303] = 144'h12d50d41f4f51da3faa506ccfe1f15d00443;
mem[304] = 144'he153ee03180002c4fc350ae20a99f23afe28;
mem[305] = 144'h0798f2b8f6471688ecbbf30c187904b7f257;
mem[306] = 144'h0cb31e1c1bf21d83eaa9003609b019a5e544;
mem[307] = 144'hf069ff8a0e03e316f04707c0f5d5ef24ed64;
mem[308] = 144'h0f5ef50dfaf2f75f0612154de119fa9bee8b;
mem[309] = 144'hf177e51e1c3ef894ead0eac317e3fa25008c;
mem[310] = 144'h0658fd57eb91e59feae2058b1b41e48613c8;
mem[311] = 144'hec2b070e18fc0c840aaa0aaaef340bd8f549;
mem[312] = 144'he6c71dd9eecffeecfb60e7871e13186412d4;
mem[313] = 144'hf8b3047602301bf314f6ee1e01eafed5f64d;
mem[314] = 144'he72fff75eb6b0d55e1e8119d1402ee601452;
mem[315] = 144'he76201d8edeef86002b2fd0f0c1af5381234;
mem[316] = 144'hfb76e30a1be217dded59eb43e9870a3ce993;
mem[317] = 144'h10d10e93f2a218d9e8be0287edaef644ff1c;
mem[318] = 144'h039cf6a603a3e56c0456ed8502ae1040fd80;
mem[319] = 144'he5a8054df914077bf9df1d08ea34e522e48f;
mem[320] = 144'hf1e913cd07e0ed2f06800c1b1e0d109413ea;
mem[321] = 144'h0af9f3a4135e1b02e28ae4791c8e1c8116a7;
mem[322] = 144'hfd67f74ffec3f5b21c3f01fdf44bf02cee5f;
mem[323] = 144'he15b077ffb280993e31af812f89807adf083;
mem[324] = 144'hf9e8f17ee2ea1a38e050e849fd3dea5ef99c;
mem[325] = 144'hf5deef3e15aee8af0e2ce7eef4dc1c20f994;
mem[326] = 144'hf2a71d3b1a68196f117ff5b71da5fdb20c3c;
mem[327] = 144'h0d571933fd96fa51fb25eb49e206f70cf1b5;
mem[328] = 144'hfe3c189be6afe140e789fddd092b1071f2f7;
mem[329] = 144'h1cf81e20e998e3260f1c090f0d491b731cbc;
mem[330] = 144'hf41b18c8f4c401cbe9d8137511f41fc71d5e;
mem[331] = 144'hf50b1e53f900fff6eeb21d54e13f0e0e056f;
mem[332] = 144'hf6b2f7131e0a16080691fa7e0ca6f1b917e6;
mem[333] = 144'hec911189fda1dffffc9cedfb0e2bdfe618b8;
mem[334] = 144'h09a809a3f7121ec5010515c311bafcb30ed9;
mem[335] = 144'h0547e5d1f7280d39153bef6cfd38eb35f80f;
mem[336] = 144'h020bf6d41b761060fb1eed9fecd3e79a06f0;
mem[337] = 144'hf2d2e0be06c0fcf2f10f0ee51b1801e80a46;
mem[338] = 144'hea170a8612de1d70165d06cdf105ee16f230;
mem[339] = 144'hf2c5f472efe5e3cf153d085de5f8e50ee043;
mem[340] = 144'he34a14681b37036709ceff7eee2eeffb1f69;
mem[341] = 144'he332fd26e67f0529ec5fe0e019deff76e984;
mem[342] = 144'hff07f8bee773198a103b107eef25ed5702b1;
mem[343] = 144'h10dfe1c21a0b0d4f161607230b53e22cee9e;
mem[344] = 144'he6fb07291e4af4c6f17ef4f3fa37f220f8a5;
mem[345] = 144'hf5411b560120f3caebc6047118d206e5f749;
mem[346] = 144'he437e9f0f977134a05301c84fc2f1f780833;
mem[347] = 144'h09be1cbf1228e0abf203f9e00c18e477f47b;
mem[348] = 144'h1aa9f82eec931afdf91af3770fd8fa1701f6;
mem[349] = 144'hefa3f119e28407c21f58ec48edcaea0e0730;
mem[350] = 144'h05b802e7006fe49c19820916e99304f015f3;
mem[351] = 144'hf85ffffaeb8b0174e72e04baf0dbe1391c50;
mem[352] = 144'h1016f5edee7f104907f1fd43f559e04df3d1;
mem[353] = 144'hf24d1893f64ef904e8c61c2cf84defa0f508;
mem[354] = 144'hfafff425fd3ef5fde8c910ebfd78ef171a7c;
mem[355] = 144'hef63f35c1be71add0c14011b1e080954e5ca;
mem[356] = 144'h1caced37101616d01d2415b8f7c5f933fd92;
mem[357] = 144'hed19fdc4151bfc64fdab10c8097e0cf618a2;
mem[358] = 144'hecd9f0b91ea7f0a6ecd80b66f7d40cbde872;
mem[359] = 144'hf16beee802f00a9ce0ff1f9f1681197c03e7;
mem[360] = 144'he88b1dcaea1ded8b0a86ecadee7dfea8187b;
mem[361] = 144'h0a8a12fafc23186f168403e11fdef6c500a0;
mem[362] = 144'he8df10900aeffc03058beadb104b152ee365;
mem[363] = 144'h11e6f5830191e0e2eae5ff46186f0030e909;
mem[364] = 144'he9d505ee09e516f012bd0858f858f50a1596;
mem[365] = 144'h0eaf05d7e18b00ef050cff29e22010bff742;
mem[366] = 144'h16ffee4ce6c31ee319cde08b04ab1c33e9ee;
mem[367] = 144'h12e30db5faf9083ff724ff90195ae6e21e68;
mem[368] = 144'he9d60fc9fb70e3a3ebc905cf034b1c5effba;
mem[369] = 144'he2301237f47cee701575012d17c5f21f01a9;
mem[370] = 144'h062618afffa0e40e0a49067107e213d9eeaa;
mem[371] = 144'hecf7e9131356eafe0625099dec2aeb480622;
mem[372] = 144'h182709e4e3de1d48ffeb0507fc3df5c51f03;
mem[373] = 144'h018418e6f22ce6bb17010e4dfab7f743f6a5;
mem[374] = 144'he656ed35ed400fc218bdf14e0a350ed3fc98;
mem[375] = 144'hf2e11c47e993e3831014f557113edff9fe00;
mem[376] = 144'hf5a6fddf0c7b178e157413c207a60fdc19e2;
mem[377] = 144'h1397ecf20fb8e24f0c6be206fb511e0eeee0;
mem[378] = 144'hf042ec51fb56f6ec119b1a381a41115ee6ea;
mem[379] = 144'h0b1c0fd70702e504ea12facceb8de5130bb3;
mem[380] = 144'hf4b0edfbe63018c8fe6b002202da194ce258;
mem[381] = 144'hf5f4eb75fa1507ba147a0d14f532f17efbd9;
mem[382] = 144'he219ef42f623e78a1b12e1a21f92f13e0810;
mem[383] = 144'h167ffd1915e9ef59f957ff3e0a0a18bbf931;
mem[384] = 144'h1d390d341526f4c1f5e1e19c0bec1486f91c;
mem[385] = 144'hf844f8351f371af0f3e2e0a704df1b0317f9;
mem[386] = 144'hf4a3f2f2fb510741e28a0e4413520cf8eff5;
mem[387] = 144'hf64a160e10c6e5a3edbf17c3ea8a07a5f32f;
mem[388] = 144'h14f804de0e38138706b2f1a4e3e21b6dffe6;
mem[389] = 144'hef35f1330184e117e91f1690151df62b04ce;
mem[390] = 144'hf39608571af7f9a7fc180746f393e502ffd8;
mem[391] = 144'h1d8a08d417cb12e81486fcb004e51a5df105;
mem[392] = 144'he5d805c0e812f80cf78315d016eef496125f;
mem[393] = 144'he4f902e21d4a1dace492080df592f3421070;
mem[394] = 144'he9590c2f05f4ee00efa6191ae8f713a0113a;
mem[395] = 144'hf2de071afc10f4f8fb4ffc35eac3fd17f0d9;
mem[396] = 144'hecea086bed0fe1d3fd430725f3cff99a16b5;
mem[397] = 144'hfe2b09ee139419f0f239e498f2e80c3c166c;
mem[398] = 144'h14c7f47606a2f0ace52fea2509fafaf506ba;
mem[399] = 144'h0ba30e05e43f1165021dea02ea58e8a2e652;
mem[400] = 144'heb8b05e2efa604450b68e880179ffd31eabf;
mem[401] = 144'h0cce08c50df30941ed060d91ec03028e0a2a;
mem[402] = 144'h1523f2e318fb03e5e961fbaf03e818340b23;
mem[403] = 144'h025df271e3f3f37d0240f52f006e1e16119f;
mem[404] = 144'hfcb60414f253fac00daaf731f74cfcf91f3b;
mem[405] = 144'h05dbe7afe64ff9110731efd11f511bf70586;
mem[406] = 144'hececf6a20ae10be2fc01fe7a1b9cf9800ccb;
mem[407] = 144'hed8900491011f29fe6950014f121f5b51bd2;
mem[408] = 144'h1a4ef8340e0ff4d11c1a0fc61971f2c5f39b;
mem[409] = 144'he50aee7ffccc00ed1b6a090aeb71ee4d12b7;
mem[410] = 144'h18941db5ecb218cb01670d29149a08b2f3ca;
mem[411] = 144'hffa20f490cc9ec74ef141b110d2d0d470d9d;
mem[412] = 144'h15baed98f643ee0ce3a71d64f929092df3aa;
mem[413] = 144'hfa6cfb3cf2a515ece7d31e1fece9eb68e510;
mem[414] = 144'h1d9106a90b01070b1369e0180d6f030c1986;
mem[415] = 144'h11f41a801f71e8461feaed1e012008e8097a;
mem[416] = 144'hf977f2b91534f1c3195002dfe7eb1fb70b6e;
mem[417] = 144'he83613b7e0c3f79014b6f4331f8b00201cc5;
mem[418] = 144'he7da1a0e17f41a03ebd30961e1960d810981;
mem[419] = 144'he7f51a2a1a070afbe39103af00870ad4091d;
mem[420] = 144'h189bf4241dba0696e4080233f81f01b30270;
mem[421] = 144'h1408ef21fce5186208dc075bf8420e5e084d;
mem[422] = 144'h1635e8aaee5fe0260bc5ecdaec071b0b01c1;
mem[423] = 144'hf85c07ca114be70c1d72e3841aa2ee7f1e02;
mem[424] = 144'h0a4713581a1c0319ea03129806831685e10d;
mem[425] = 144'he3b30bc01e0b1a6c036102eaf82efdefe4fb;
mem[426] = 144'he74ee48ef7ebe2db0374fce2f3ece90e1960;
mem[427] = 144'h08e20210fc35f5a217ccf3b2fc680e591c7e;
mem[428] = 144'hfdc7e4791007ecc8f3fbf9061ca80d141039;
mem[429] = 144'h02371e3efcdde8b502e8fbedeefdfacfea31;
mem[430] = 144'h04bf0592fcc7f227e142ea8a0471e76c11f9;
mem[431] = 144'hf92b06c001c609010537fe1101030949f897;
mem[432] = 144'h02aafb68f1a206a0ffca0a4ee934f5c717ed;
mem[433] = 144'he4c0e43808c818a306c2f4ed191efa3b0783;
mem[434] = 144'hf013ff8b0885ecdf094ceb4f12c90a4f0d08;
mem[435] = 144'hec56e73f09f5ed16fb96e1d5e34bf53ceb7d;
mem[436] = 144'h16a3e953e98f017aebad1c0cf3480013e881;
mem[437] = 144'hf8bbf070f347f2940ff8e31cff1015020694;
mem[438] = 144'h0caeeddfe9a015c8e72505aa0d98fbefee64;
mem[439] = 144'h0abcffcfef3d1872fad30356158af75eedad;
mem[440] = 144'h0560fa720f2bed4d143a1b9a0a770408ea7a;
mem[441] = 144'hf7bf1730fffd04ab020f16260dba0cc01b6f;
mem[442] = 144'h1ba919faf91af48ff599e00bf1621a5414c6;
mem[443] = 144'hfca40f9512a5f29df29f03b21fb6f08aed95;
mem[444] = 144'h1d6a0aa9eb641d06e130e825076ae5f9f678;
mem[445] = 144'h1beffb02f1e6fc74e3990899ff79190118f3;
mem[446] = 144'he84bfd32036df2f719c81faa1c421f09e06d;
mem[447] = 144'h0fcee47b00611fd81fe5f9d51442e9a10c17;
mem[448] = 144'he9faeeebf882e801eb8a1f06e547f2b01fae;
mem[449] = 144'he5bf17cae73208540e56fd2be1590903e2b4;
mem[450] = 144'h1c02ed42f2b4126916d11818f17afc221593;
mem[451] = 144'hff4507491cab1e63ec35ee23f77dfd4ef222;
mem[452] = 144'h0975e855063906ee1831f2221ac713dcf5b5;
mem[453] = 144'h121ae50807170b8bf00de7370779ff3b0d48;
mem[454] = 144'hf63806c80de812ab03721708e6a5ef30fe7b;
mem[455] = 144'hf7f20715e87a0519024dfca01b8a051aea0b;
mem[456] = 144'he9e2f128eeaee6870cc21335fc7ef817f043;
mem[457] = 144'h08310040ed8e0e25f4c5131e07c3e5ba12bb;
mem[458] = 144'h15cee5940097e95518a5e30d14dbf142eca0;
mem[459] = 144'h07dfe2aced6d12b8e7c3e501f93102ec1159;
mem[460] = 144'he0d6194e0907f82efa8d1471144cf624e02c;
mem[461] = 144'h1de0ee5d1e7af57be1e6f6430a8ef62b0a25;
mem[462] = 144'h11ccf111fef614fc16c1feb2eb97f90213be;
mem[463] = 144'h0243fc92eea809fd050ffb73f2e013ebf722;
mem[464] = 144'h1b4df302fc05f5c4e82ef0ef02eeeaf8f67e;
mem[465] = 144'h07f11ccb16ea138df513115dfb150d3ff19b;
mem[466] = 144'h09efe1a9f2aff64616a0f01d14aa04070e8a;
mem[467] = 144'hfa0df22c02e8e289f4fb1247056de19ae8b4;
mem[468] = 144'h006f15eefdc5eb3d124808f3fe8d13820ea8;
mem[469] = 144'h0dc30ad1f66a0f1b0337f61ffa1d04450dc9;
mem[470] = 144'h0a46fc11e655f1971e130f55f3fdee86e2de;
mem[471] = 144'h0bb8e6c01239080cfdd3ebd718b9fc0afcdf;
mem[472] = 144'h05b1f056edc0f183092c0e7ae94ce5b8fe28;
mem[473] = 144'h1554fea9006919d10ed31821f330e1f90503;
mem[474] = 144'hfd9500681459068bec13eda6ef201f5c182a;
mem[475] = 144'hf2330743142a1da014c01cc615e51e9f01a9;
mem[476] = 144'he8491f65eb791ae709d6f71703c30c791b66;
mem[477] = 144'h09a0138bf2f81fbaf215e078eff01effeed9;
mem[478] = 144'h1e96f146e1430909eb8bfcb402450049e593;
mem[479] = 144'h1425fa2b0e1afb131bac1080e0ff0cd4e973;
mem[480] = 144'hec6df98ae8eb040909b9e64eed4cebed03d0;
mem[481] = 144'h0782e85d09020fb3e1ca0dc0155cef3be41a;
mem[482] = 144'h102eeae1efca1df2ffb7f6d70c0f1f59e13c;
mem[483] = 144'h0f080083f388ff771c02f29c1fa80178040e;
mem[484] = 144'he4ddfe60fa5301281c14e26aeb8be78afa9a;
mem[485] = 144'h1ff90176069019481baffe4907ef0e56fa0d;
mem[486] = 144'hf88ffe7d039d164e06a6164c128af1641432;
mem[487] = 144'h1e68ef3718a2e737f21de77310e204b0efe5;
mem[488] = 144'h084511970da5f8be048e0838050afe27f841;
mem[489] = 144'hf88ce6f2e2eb1219f3a10db00bc4012be439;
mem[490] = 144'hec4af6a8e52c1b1a05d0fe7fed7dfd27ef78;
mem[491] = 144'hfc54e66cf786f76ae9a0e7d7fc86f6eff453;
mem[492] = 144'h1aa40ae606f60fd5ed62f045f1f1fccc1d77;
mem[493] = 144'h125b078013d31ef3080517fce8fffe3d12ad;
mem[494] = 144'h05581f8af0b0ec37fa0108c81419136c1d4b;
mem[495] = 144'he8b003cd10ba0e13ef75fa5e1df90edf0262;
mem[496] = 144'hfffc1c1bf390f4eb19581643eeda07e3e2ec;
mem[497] = 144'hf59c0710e690fda61640088509ac1bc30b4f;
mem[498] = 144'h13e5f3590d14158111f9f36a06a61d44055c;
mem[499] = 144'hf332027de5aa0905163be3a9fbd91f4fe93b;
mem[500] = 144'hf732eed4185affccf3371076f30307931b2f;
mem[501] = 144'he14c0bc116890e0d1cd1e51706d80aaaebd9;
mem[502] = 144'h02db18c301adf35109da00efe93f13d9ecca;
mem[503] = 144'h0acfe119f679ef230fb3e8ac06e602c8f0f1;
mem[504] = 144'hf1fb0d3d12560d1de014e1ca1f720affe237;
mem[505] = 144'h00af15670f890574ed87eab6f09f18730962;
mem[506] = 144'hf025eeceed0ff9ffe8aae312131f08ab13d6;
mem[507] = 144'hf8bff03102431791f149f816e292155e1601;
mem[508] = 144'hec531ba2101ff8baea6d12d513de06c20907;
mem[509] = 144'he325e0e7e51bfae00b87e0c502ccfdd90f09;
mem[510] = 144'h13640956f3f20519e3c7fec312f51db5e0b4;
mem[511] = 144'h16fe1130ed8b1b92084c0575fb0c0c5dfd4b;
mem[512] = 144'heba30859115e00e416cee165040b0a1efc8c;
mem[513] = 144'h0aace95cf31ff5080a8fea70fae0ef02095e;
mem[514] = 144'he3181d8711ad0d84f1831deef8c0f5861af1;
mem[515] = 144'h13a7e354faf3f9ebf06f0cba0c890e4a16c0;
mem[516] = 144'heeca11fdee64162816dcebfe15131174e480;
mem[517] = 144'h0a28ff5816a6084006770ba3137aefbae16b;
mem[518] = 144'he8ece0e0ed7ce90d0ad0f5d5f41cfc700148;
mem[519] = 144'h0c98153002231f06e2f91cc00fc408931f27;
mem[520] = 144'he9effbd2f9cefb14166df8e6f725fa001f87;
mem[521] = 144'hf1920baae0b01294e9b51a6be2cae6c1eb1a;
mem[522] = 144'h148111a2108c1db30ea20c93f37e0a361b47;
mem[523] = 144'h19c60ff5ebceede9fbae1aebf226e60505e9;
mem[524] = 144'hfc1b0427ef741cb00cdef44be9abed6bf8ff;
mem[525] = 144'h0b6510d91985164c086aec57e66415ce020a;
mem[526] = 144'hefdafeb81afa159ce608e853110b046cee8a;
mem[527] = 144'h044600be087a1c0ae8321188e08af078e31a;
mem[528] = 144'hf9a61a06e20e015af6d51ad9119d17841e9f;
mem[529] = 144'hf7871a3c10fe0172e1aa050c1004f0a61b71;
mem[530] = 144'hfa8a122714acedbf1de9ec4fe431e9f2e5dc;
mem[531] = 144'h1a79fbf8f785e3a7f82408dae10df967e1f2;
mem[532] = 144'h170d0bad02c004a91456009e078ff23bf848;
mem[533] = 144'h021af21102f50b5c13e6019e05cef32dfa13;
mem[534] = 144'h0a6f05030aaf0c9ffbc8eb99110c1a480eae;
mem[535] = 144'hefd5ff92f9b216a401320311f312190303c3;
mem[536] = 144'h017df76013c205f61033ea6401870995e6f3;
mem[537] = 144'hf935e4e2041a0fe0e6851148ee1f10abeb37;
mem[538] = 144'hfae603f11813fabdf0811369f817e372eada;
mem[539] = 144'h18dde97c1194e4221d891c14fe011fd5e720;
mem[540] = 144'hf50d0c73e5af013a1efceb6b180c025213fe;
mem[541] = 144'hed3deff5f00f1c15183603cbef990e47e5f6;
mem[542] = 144'he086083af19fe9a2024501d0e634e72102b5;
mem[543] = 144'he54a003cffa0ed41efedf5ae1dc51dfdf906;
mem[544] = 144'h0b691499f6830c931626ff08e7e714d8edad;
mem[545] = 144'h1ec40a78f3e6fc50ff52ed11e45b0387ef6f;
mem[546] = 144'h0e6e0b171398e0fd1f65e6431fe9fab1037e;
mem[547] = 144'h10f8ee00169008570ef20974e9c305cf166c;
mem[548] = 144'h089aea511ca6eb44152505e40a78f139042c;
mem[549] = 144'h1d43018a08e00ed6f3f70104f176febc176a;
mem[550] = 144'hfe16e441fcf0ed4100a4e53df32dfc7fe3ba;
mem[551] = 144'h17d700bfe63f1a32ea86e5c30e2902aa1641;
mem[552] = 144'hf09917bae3ebf3e4e6eff2def67f1dfd1509;
mem[553] = 144'h12d5ed57efe1f41ceb8bf57107461624fc37;
mem[554] = 144'hf2d2f29518c21d310646fe07e144e2bff81e;
mem[555] = 144'he723f2490def096712ee0da5fada0f6c1138;
mem[556] = 144'h1074feba1551e88d0961ef31f173f9beed5c;
mem[557] = 144'hf8b40566f02dfcdfef90f376e4941b4fe59e;
mem[558] = 144'h1bb71655101e11e60dc4fac815c70ec8096d;
mem[559] = 144'hff90192cfe8efb49f08200761919f05517ce;
mem[560] = 144'he406f05e0e66ebae1933edc6edefe1f3fbef;
mem[561] = 144'h00bfe590114217e504fe1bb6f6bdf147f6b3;
mem[562] = 144'he8e615cef03eed71e5680c680a4f037d1b93;
mem[563] = 144'hf5641ac61ef9edbc1210187d199204afeee6;
mem[564] = 144'h0ed0e90909d0e84dfbdeef4d0770fdd5106c;
mem[565] = 144'h0c811b33f4391984f16d1c31fdbc1d4d1802;
mem[566] = 144'hfc11f2b8ff62ebfdeeb8fda308cdfa81faf2;
mem[567] = 144'h11b5ee7d12af0ac9148e14e719b41e81f4dd;
mem[568] = 144'he5190fcfebad0e9319040adce0e0eaef1c29;
mem[569] = 144'he66b0eb6fc28002315ae1909f08fe5bfed3a;
mem[570] = 144'h187de5cc1c7ffd0de30ef9790610f1c20989;
mem[571] = 144'he1a9e29e1629e33506d5ff29ed261d33efc3;
mem[572] = 144'hec5beb09025df96808f21b9b1ebef4191226;
mem[573] = 144'h1693f9b00bd5e919ecf9f1460759024c0069;
mem[574] = 144'hf8b6ef920a730b33ed6f1d7a043a152aec4d;
mem[575] = 144'h1e2bf06211cb00e8ea271bb71c36fe07ec36;
mem[576] = 144'h1fbdf8b1fa25e984e532ff001556efb6035e;
mem[577] = 144'hf694e4ba1b31e07805e405531d49ea29f4e0;
mem[578] = 144'h087cfaef133b0256f51ae625eeabe1e8ecc4;
mem[579] = 144'h0e0a0c41e373084de0bfea80e2f8007e1051;
mem[580] = 144'hea020acde22f0a100299ff18f0b9f7c30ef4;
mem[581] = 144'hfdec1034e4ed1b89fb72e86ffbad09641386;
mem[582] = 144'h11e1ff2afde7f7de034ae5d90e8405c5e518;
mem[583] = 144'he8f8ebadefe611f3110dfe78e2d5f91fef02;
mem[584] = 144'he2ebf2caf196f609f6db1857fbb6e81a1569;
mem[585] = 144'he9e9eaf914070f6cf5a015e6f5a1f4891478;
mem[586] = 144'h179e018e1356e4f3e6da0629019ce4c1fe58;
mem[587] = 144'h0abb0a41f98109b505f2f6b715141ed9fc74;
mem[588] = 144'h0e00f808e4ca179015be08c0086df7dce766;
mem[589] = 144'hf24fea02046810adfd7ff570e50e114fe6ec;
mem[590] = 144'h05d0e8e2fe8dfa3a0251ec59ef9a1b1e081f;
mem[591] = 144'he256167a1b1002df0cc4e5e9f2cb1a10097c;
mem[592] = 144'hf312e80614d80dcc0dfbe660f5d21272ee58;
mem[593] = 144'h0c1b19b11b781bdaf1f4057f1c26f0a0029c;
mem[594] = 144'hefd10d0f085be71cf12eecd1e5eb178701b9;
mem[595] = 144'he22ae771f6f3f944ee330aade1e5e956e3a2;
mem[596] = 144'h1cc70a29f8e3eda41a781aeb17d7feacf866;
mem[597] = 144'hf30a0067e080fbaf103a09caf7060c0a0367;
mem[598] = 144'he73feb11118d0e2205d405bb0d94fc6500f7;
mem[599] = 144'hf0621b1dfda01afce9f11a32f62af59e0e6b;
mem[600] = 144'he4e7f1431ced1ebce9ece477eff91ae4ea87;
mem[601] = 144'he367f34c160102b60ff8ecedfda2eadb1158;
mem[602] = 144'h145df62e18720e04ec8b0717e1410885e6cf;
mem[603] = 144'he84200df074e0916090d1b251435f758f4af;
mem[604] = 144'hee751263fea9f3f610edfc84ed92e30ff14c;
mem[605] = 144'h01dd0d04edda1030102915bd01b811e81676;
mem[606] = 144'hff48f25af5abfe7c0c0517d41ceefcd80271;
mem[607] = 144'h15c0050df36204281a6602bd008a04cd0eb5;
mem[608] = 144'h0b5f13f6e15205b9f208e4b3f160f98de700;
mem[609] = 144'h082eecad0329ec4be8310b17fc6116671089;
mem[610] = 144'h15c0fecdeeea1689edea06d9ef6a1937e819;
mem[611] = 144'h0766f7031fe512f3e44af88604c3f2a00d49;
mem[612] = 144'hf9a0093417eefc820641f734e058fc0c19e6;
mem[613] = 144'hfae818a4093ef73bfd5215da1a441b9f0b85;
mem[614] = 144'h0c26ffd4f73ffac113fe15c80a88e4b70433;
mem[615] = 144'h038a1ca0f24aec831672ec79ef11ffc7e949;
mem[616] = 144'hfeaefe67ea8cfa4b127ce88d0a260de5ec3f;
mem[617] = 144'hfc4418371ddc0cc21a3e110bf471163afe0b;
mem[618] = 144'he2be1090e978ed0c02f8e905f8a3f6220c6a;
mem[619] = 144'hf9bc0287fd7209a013bc0626f9ccf1c7e056;
mem[620] = 144'h0826ef4f12350d03f5400ff8018be727057b;
mem[621] = 144'hf83e14b91ace1583ea95f705ff8310310f63;
mem[622] = 144'hee69082de21606101b4f0f2d072c15991cb7;
mem[623] = 144'h12a9063b096de600f56c179c192d0b240fea;
mem[624] = 144'h16bd1d68112ce93a1d0cf32018fbe6340add;
mem[625] = 144'h1fc6ee1bf0a219c3eb8713ede51ee8101469;
mem[626] = 144'h158e1489f85f1a5211210d7519c7ffdc0ff7;
mem[627] = 144'he72ff397fa9218430d2a0c5ef5cb0017ebcb;
mem[628] = 144'h0721ebf4f8da0fb1e071e411f760f056ec5a;
mem[629] = 144'hf9631addff531cd11f76f618f6421ffe0b7c;
mem[630] = 144'he3f107e80e4df32e142de299f60ffc9bf2cd;
mem[631] = 144'h00ae0369e6540e1bf2dafbdce49a11480613;
mem[632] = 144'h0286ebfff717fec702230385f9980a9bf732;
mem[633] = 144'h1f1111da024d0b240136025ef78aff1f1b31;
mem[634] = 144'h0bc1e4e21e240f8d0293112af62a0446f29c;
mem[635] = 144'h0b9805f8f2ea03711ae2f276ed5f1074e40e;
mem[636] = 144'h0330110ee3910700127df15b130fe169ff3f;
mem[637] = 144'h1cbde64ce9790f5b0c9fe228e99607711d94;
mem[638] = 144'h0c65ed05059b18ef187c04b70e27096dee15;
mem[639] = 144'hf5360283e5fc0f37e55b029df66205101d8c;
mem[640] = 144'hec0dffa410a103d0fddff6b21963f69e0d31;
mem[641] = 144'h1e6b0b7c1780fd9c1c1ee2c3f7a311a306c9;
mem[642] = 144'hfcfdfbf6fcf3f521f76418f7ede8ed61f415;
mem[643] = 144'he33bf353f85811e7180ff376ee07e90b1fa5;
mem[644] = 144'h131a149d0fcd0a98f16e06d105e3e90818fb;
mem[645] = 144'he69dfd15e3141d4715d3e438026ffab413bc;
mem[646] = 144'h053b0ed9ea0e0b4bedc2f8a10fd51a05177a;
mem[647] = 144'h1e7107cf0521ed4b0e2e0c0cfcaf056e0bae;
mem[648] = 144'h172bfd9cf50808c9f35a197d1a71151e0afd;
mem[649] = 144'he64eff5ff0c310a3fb7df8e1fa900cc310cd;
mem[650] = 144'h156e0251faf6065fff3d129be77ae0330a22;
mem[651] = 144'h00d90badee2cecc619380609e7b8ff0be399;
mem[652] = 144'he6dae47102cf0a95f864ff970974f7201b1d;
mem[653] = 144'hf6c4eefcf5a8ec8802fee91bf3c4157d0254;
mem[654] = 144'h10be0a14e37f022509391220165bf65ef76e;
mem[655] = 144'h10801736e9be0bf805f7ff68ea5b0b7c1457;
mem[656] = 144'h16f6e0fdf4c8f2531c3de74d176811a0ff01;
mem[657] = 144'h10dd02440f4b18fdf627191ee318e19e00d2;
mem[658] = 144'hf944170affe4fe07e9d5067ffeb10e2febef;
mem[659] = 144'he38903efe6b20cf6f1c2099419dbfa030112;
mem[660] = 144'h0bee07480f6ef329e8cceb241b31f109f086;
mem[661] = 144'hfe9af46f032ce45af43ce081ed2c10c0e83e;
mem[662] = 144'hf7bf1f4bffecf53d0ce001ea11d3001b0f19;
mem[663] = 144'h11d007e6e08c0d97000b187ee4780bbf1c63;
mem[664] = 144'hf2ab1b8314b0116ffa6fe0b5fa5c06f61ba1;
mem[665] = 144'h1450e452e0ea08f1ee83e6e01d980049030f;
mem[666] = 144'hf0c20b8fea4be837e95ee266016de4ba1550;
mem[667] = 144'h026ff4b4141c12b2eb1d03d7fd4516bce6ac;
mem[668] = 144'h091bf0affb38f6fe1ad709ff0fcb0c8a0252;
mem[669] = 144'hee1b098c15ff0e7fefb2f327eb83f1591937;
mem[670] = 144'hf553fa0eeed9e76f15f91524e16616b8f907;
mem[671] = 144'h16fdf59d15ee132fe7041c34fd0be2e4f7d2;
mem[672] = 144'h0cc218ccf67f0bf9fb4001da01c009c6f5fa;
mem[673] = 144'h183bfa97ee4ae768ef8fe621f97407941fe1;
mem[674] = 144'h1d8be0920299e02fea9017321a310cc81ebf;
mem[675] = 144'he1ae12f305bcfaec0c57f7030bb805f50271;
mem[676] = 144'he0011baaeeb511720d5b0867fd50f64efa79;
mem[677] = 144'h11acf58ef5f1f5e2eb6ee06fffe0fc9eeadd;
mem[678] = 144'hf6fcf9bbec951cae1856097e0b56eaa20a75;
mem[679] = 144'hef8cf2b5ef320ed20f80fdce19dce89c129f;
mem[680] = 144'he0430175e9e7f0a00edeff9bfad7f24be9e5;
mem[681] = 144'h0838fe5f000d027ff823ebdb05fef2cded9f;
mem[682] = 144'he48c10a9e9aae5d3f4bb102718ac100d071a;
mem[683] = 144'h108117d6e6a6e52aea4f00041d07f240f771;
mem[684] = 144'h1b8be802e9aafe44166e1543e3100e76f376;
mem[685] = 144'hf1b20d42f5050414f2b1f7a61c28fdef17e6;
mem[686] = 144'h091d1631ff53e0defd2408e4e51d0bfeea89;
mem[687] = 144'h058fe381e8ea11e900e80d20f0dfe9b20cc3;
mem[688] = 144'he09c1dcc04d9098511460106fd8be1291d4b;
mem[689] = 144'h1f36e5200f6604b7fd3d1ae0fd98f163fa9f;
mem[690] = 144'he0831fbdf5ebf3af19210b3eec65fd790d9a;
mem[691] = 144'h1d24fe11e95a0933e8e51a6cf7c613cbf15b;
mem[692] = 144'h002b0a551b20f6bfe2a8f6d6fb26f029e036;
mem[693] = 144'hfe3eefe0e09ee05c164ef2abea710ac40c9c;
mem[694] = 144'h0dd01872ebb2e754f0f9e6feebd4ec481d8e;
mem[695] = 144'he59619491f2dfbe6ec99e53bfcc81e91e8f8;
mem[696] = 144'h02c7056b019beb4bf81ffd28e95de2d81b94;
mem[697] = 144'hff5906e9ef5806b41fa4e2fefcad07e50356;
mem[698] = 144'h0670fada02dc0ab9e25bf8a31e3be317e40f;
mem[699] = 144'h162fe06ce5c9eb00e1fdfd87102ee9d7dff3;
mem[700] = 144'h0059f7b11e8e0312f9711406ee67eff502b5;
mem[701] = 144'h0d5ef243fe10f7f11457ed3b1549f56803a5;
mem[702] = 144'h08a510f3136cfcadf3710168144f197bfde6;
mem[703] = 144'h0806f1f61c8302fce480eeac1e3ce1f0131a;
mem[704] = 144'h1f8a07d60829e73a0e7ce81702fee99210a2;
mem[705] = 144'h15c1ff0ffab0ff62fcdc1bac0742e1aef6f2;
mem[706] = 144'hf980f197f2a1ff011c85123afcaceae914c9;
mem[707] = 144'h019d129ff818e502f7fcf8e1f9abfe1af835;
mem[708] = 144'h1f14eff3eb03e5c5fbf40c3b09ebe12202ef;
mem[709] = 144'hf46beefa08f8f9091697edd9016ce5fff630;
mem[710] = 144'h0caaec140b4e1a6a15e8107ff38601c818cb;
mem[711] = 144'h136ae1190f7c171513c60b9001c7158c103c;
mem[712] = 144'h07981786f8481e4ef51a169dfff6171c13db;
mem[713] = 144'hfda0ff8bfbab130df25afd30f180089fe766;
mem[714] = 144'he22befceebdcfb5ee44afab90ed100e9042c;
mem[715] = 144'h1a37146e0871046ff57100cd1f5be0b70f88;
mem[716] = 144'hfd61143e16bbf607f9bcfeb0e2781521dfa1;
mem[717] = 144'hfc9df14607ca1a6df8f41bf208fc0095fc5c;
mem[718] = 144'he59b1f3ee7be183aee6e061b0a20e703fb57;
mem[719] = 144'hea9ff974f71afe9414cbe42ef525150d0f8b;
mem[720] = 144'hf150fd0ce0daf5fa043613c113920e570e91;
mem[721] = 144'h1ccaf81af3520409ee9ef099f6c9fa0fec1e;
mem[722] = 144'hff3fe2300d27f0d7012a026f078c12de0bd9;
mem[723] = 144'h106bfad21bf2f86215800b68ed230b2c00cc;
mem[724] = 144'he073e2fd15230e8a0b8be38610e9fcd9f615;
mem[725] = 144'hf8d6f78c035f06bbe796f3950dc20c2b0892;
mem[726] = 144'h13030aa219591b531388f938f41a1a851b7a;
mem[727] = 144'h0d22eb0ee5da11e8169de5dd1e4ae29bfa24;
mem[728] = 144'hf7f1fc4a1c531388eae40957f8bbe422eb1e;
mem[729] = 144'h027b1504e105079be8971be31073116f1cea;
mem[730] = 144'h0264ec8cf331f075e2a9f77c01f9eb511d37;
mem[731] = 144'hff7306421163f1120fe1fe28e0eb0698fb76;
mem[732] = 144'heaf7f17416110121ea220f1ee6f8005008e6;
mem[733] = 144'h0ed3f560f805eef0f4891dba0bc71a40f8e3;
mem[734] = 144'hf17d161b085018370ce3f41308010c9e01ef;
mem[735] = 144'h043d1dcc0cedf8641eb807be1cf00a63f297;
mem[736] = 144'h14b002a615dcfad80c130ca6f1b9f57008a6;
mem[737] = 144'hf675f03ce5f81fbde450fbe312cb0d290c38;
mem[738] = 144'h078fe9bc1bc60bb8e12de049060818dd0c1f;
mem[739] = 144'h05bf0f540cd3fc030c87102cef36107600fc;
mem[740] = 144'he29fe261fa4b0ddb0350f4ecf84c19e50951;
mem[741] = 144'h0d34f220fa8be9651075061af307f223150a;
mem[742] = 144'h0570ff53068be0e1f76ae2431fe3e2490d9d;
mem[743] = 144'h1b3d02b4e465ec39e9f6e399131de497f732;
mem[744] = 144'hfde1f4a91ce3f4b6f811f3aff357ff3104db;
mem[745] = 144'hf74fe31b06cce38900b5020df99e08f110cc;
mem[746] = 144'hee47f4650eb5f940040bf4601ffc10d4f5ca;
mem[747] = 144'h17821ef71cc2f2c0e23a040b01d30b9bee83;
mem[748] = 144'h0c05e55f15fb1c3ce3520a18f8d6fe060c03;
mem[749] = 144'he568fe3d0faa1b8f00df183b08e002d81e84;
mem[750] = 144'he7c51a430368e34c0be516eef215ed2f014f;
mem[751] = 144'he876e805fc5f0fa4f76fef250a5902c5fb23;
mem[752] = 144'h0cc0f7e3e1251920f5fde849e86ef9a6fcab;
mem[753] = 144'h02320beb128419b7004d03fc1f991b9f10b3;
mem[754] = 144'he47bfeb206071a51fad6ecb60a9ee91f01fa;
mem[755] = 144'h0f4af6e2ef8cfa0b0c79ecc31899eba8fe03;
mem[756] = 144'he69e0df8114de530eb630738fd0f0a0d1ba9;
mem[757] = 144'h196f1f151381f9ffe8e7041405ecef00f07f;
mem[758] = 144'hfd1ffe13f0a2e2270edae401124aea7ce555;
mem[759] = 144'hf9c2e6bd12c7fb750c7e1f370191e564198f;
mem[760] = 144'h145810551fa3f55005b8e3b111c40893e456;
mem[761] = 144'h0bb6f360f186f5ed0ef4e1aef7390c7ffb65;
mem[762] = 144'h0b35f9821d81f3ce0215fcc7f624062014a2;
mem[763] = 144'he8fbf2311960f23ef64c0a5cfe631f730a7c;
mem[764] = 144'hf884e2641332ef4401a41583e1a9eb1bfb6e;
mem[765] = 144'h15daf1181a01059c05ca0a7ee605f8a3ffdb;
mem[766] = 144'h1343fee5187d1168e193efd719761210f614;
mem[767] = 144'h17920eb208f4e19901d7feda1a48e4401068;
mem[768] = 144'h13c618bfeaf5f3100a94fa6c107e0ed4fece;
mem[769] = 144'hf80de9d717fe02741015ff79195be3d2f8e9;
mem[770] = 144'he92218e305f50483e7d0fc14f1221c24ec16;
mem[771] = 144'hf4711cca0f7ff186169d0b6a1af607a8e9de;
mem[772] = 144'h069eef94f5c30f23e57a1ee70934e92e059d;
mem[773] = 144'h1054ff7fea26e4d506daedf41605f097177a;
mem[774] = 144'hec17f8a2054602020468e0a40cd4e9f9f048;
mem[775] = 144'hf055e280e049e4e207e9eef7f474f485fd45;
mem[776] = 144'he55315bef823ed35f5fee7f0e7fa0dfa1e44;
mem[777] = 144'h1bcce0861a2801d5f43f080efa8dea7100fb;
mem[778] = 144'he137f562086cf59b058de08bf7611955e4eb;
mem[779] = 144'hf0a00430050df62c1192fda51ccf13910f27;
mem[780] = 144'h0482f892fdd10cb5e59f049cf25ee9bdf3b6;
mem[781] = 144'hf24705791ed4004bec58e14ee89e1e4cff44;
mem[782] = 144'h0b0cfe7c1f61159509f605f003ce032cf6fe;
mem[783] = 144'hf1c81e9c0c48f0be01c4e2d0e819fa3c0ec3;
mem[784] = 144'hf1d61d32e6af02daf4960bf8e77df9ede550;
mem[785] = 144'h086f1b21e6f5e658011a0acee817e497e19e;
mem[786] = 144'h09dff2240f47f0fa1ceb03bbfb21e004ff8e;
mem[787] = 144'h16481002f4e8eecef2db12a012071146edc5;
mem[788] = 144'he2f5e953190ce55cebf4fd190f0df08bf0ae;
mem[789] = 144'he8af0c361024076812bcf8ff19b41e0b1cdf;
mem[790] = 144'hea9ae970fe870f36f44904dc1563ff42f647;
mem[791] = 144'h0f5bf4a6edc3eb0be00813fc15a5ea5aeaaf;
mem[792] = 144'he44f0500f8630b95f1721c430279f68beeee;
mem[793] = 144'hff6514f616e9f574e40e09bf02b01daff186;
mem[794] = 144'h1628f057ed7a014cefc7f955e0b414900405;
mem[795] = 144'h0c5fe40e0874ed60ff32f7c608c3f2bdecb0;
mem[796] = 144'hee350d02ff9705a1157fe3c0197cfdfdfed8;
mem[797] = 144'he06b195b174ef9c50cfdf1d2f477e0691653;
mem[798] = 144'hebfcf734e2361047181df2c21ed0ec2e0a68;
mem[799] = 144'heb3e0713ed2e1194eeb81805f4270af80417;
mem[800] = 144'he570166afee0f9ade638ff45113e133bffd4;
mem[801] = 144'h1fe407baf286fb45f5b90cd0fd23ef31ff20;
mem[802] = 144'hedf9122ff7d91b6af14bf8a61328fc1503cf;
mem[803] = 144'hff98e141f7ad0f3a09a90e7aef7cfaf3094a;
mem[804] = 144'hfb00e2d016bf1911f79af037089112a41999;
mem[805] = 144'he783e9e1ff02f4e1ed4bf59a11e6124afd19;
mem[806] = 144'h1828144c17880c62f4e810b9f767f863195e;
mem[807] = 144'hf9f51ad6f146053dffb2e912e3e8e35ef5ba;
mem[808] = 144'h14300aa20aabec7cf00717b916830da218a5;
mem[809] = 144'h05021adefb6404bf177b062a0f000a5ae027;
mem[810] = 144'hedd6059de860ee9d102800e8e07d0ac91cad;
mem[811] = 144'h1f6df3f7ef4cf40be600eadd1a2cf78be807;
mem[812] = 144'h02001622ea9e0122e98512c60668f30a19a2;
mem[813] = 144'h1073190719a20a7d1c00e2a3ee8eef7e07f3;
mem[814] = 144'he3971a85fae2faae1b52f23ffda0e7051de4;
mem[815] = 144'hfaf5ed43e96df0d41ac70f1d0f0b1bb0f0f8;
mem[816] = 144'he16f1455f74b0ecde3f8081c1a82f063edae;
mem[817] = 144'h040812900f71eafe1b3f1a37e1afe7d3e372;
mem[818] = 144'he7a0eae8fd02e41d193209661babe0b71503;
mem[819] = 144'he7591055ff8a1848f31deb36055afc1806cb;
mem[820] = 144'hf6c613c4e87118d61b97e262121c0e8de11b;
mem[821] = 144'he61bfc5ffae7e573e20d0fbcedff0d31f4e0;
mem[822] = 144'hfb64e70f0b4002f7f96ce592151a11580e03;
mem[823] = 144'h02830d1b0d08f4f0fa83126fed231ed4e33a;
mem[824] = 144'hf012fd26e80ff1bf16d4faf6f7b901f109a3;
mem[825] = 144'hf2cf1c9bedf7eeeb0a2a006e1ea9ef131476;
mem[826] = 144'h10d10995e25a1fba118914dbed5607c60003;
mem[827] = 144'he250e3d3fd8ced4ee6811afbf746f4611f87;
mem[828] = 144'hebc313fce877f22cf729edf2e3a004c2e696;
mem[829] = 144'hf4f3f2d9e42aefc018141fff178cea471f2b;
mem[830] = 144'h189ee3d7f82decde10fce61112a5036efa73;
mem[831] = 144'h031afc66f936e2b5edbc16a4190df6da0c1d;
mem[832] = 144'hece405a6f7820faefcf0128e1e61f13903f2;
mem[833] = 144'he2afe42ef4d11775e48d007a1e7ae4b5fd8d;
mem[834] = 144'he2c30ece009a0815194b057cfe10ef02ecfc;
mem[835] = 144'h13fc1a5becd711701c76e69becebff48ebac;
mem[836] = 144'h0ca715ce0bac04700c960425e23514aeee96;
mem[837] = 144'hf170ea460b991031136af79e088a1edfea1b;
mem[838] = 144'hfa5f143206e1f4cee67be4071111e905f0b3;
mem[839] = 144'hea2908e2139814cfe3820262f2300c86e5fe;
mem[840] = 144'heed7e7c2faab08b40218e263f68dec13f997;
mem[841] = 144'h0999f4270279e9f4e94fe45b0f66edaa1349;
mem[842] = 144'hef2ffe58f671e3e702e9efe510c21f46f610;
mem[843] = 144'he5c1ed68f4cef86f0d5eecb31f52eb9beb1b;
mem[844] = 144'hf60de1d1166a0b8ff14f1c080cbd1d8b00d5;
mem[845] = 144'he025eea214ebf64916be0f29edfe011ce8fb;
mem[846] = 144'he53b1f8af850f756ef71ee5ff5b50504182d;
mem[847] = 144'h1728e35ee17ff7bbf824e08a067bfc40ed38;
mem[848] = 144'hf4e8ee61ff16e25908bf1c6603f8e8f4ef3f;
mem[849] = 144'h11c9ea3af9581bafe2c1f2c80c18eb7d0e5b;
mem[850] = 144'hea98efc91b701cb111a2110cf39a0d3f01c7;
mem[851] = 144'h0aadf642f267e24b11f81453e822ede11788;
mem[852] = 144'hf73beeb0e9931636eaa5e2ede6751bec0de1;
mem[853] = 144'he332f9a91f8f0fb8e279fb160d9c0c3c13d8;
mem[854] = 144'h000614811856050cf15c08f8096d0ae7e835;
mem[855] = 144'h1e0ee5800a310f7c0462ef140ee90d7aea74;
mem[856] = 144'hf7a9feb5e813e68009e211cc1dc5e7b1fa94;
mem[857] = 144'h193a12450bd510ac0993e93f1e841eb30e3b;
mem[858] = 144'he49cf343ebd5f69f15aee08312bb0506004a;
mem[859] = 144'he1a808721474066ae62df19806d0f4d4ed9c;
mem[860] = 144'h1eec08c0fe9a08d5f4cbe253e8d21be9e6b8;
mem[861] = 144'hea5f191aecc60732ec1efa82eed0129be070;
mem[862] = 144'hf243f8780521f5911fdf1d14eda5f151f022;
mem[863] = 144'hfbd607cbee5202bd11070e4bea920fcc1615;
mem[864] = 144'hfbb0ee02faec07c8e2021352f14a04acf8ca;
mem[865] = 144'he9281afd021910f1e37402aae8a317e208b4;
mem[866] = 144'h00b6e53dfcf3011a1a2aeb2efc1f0c6d13da;
mem[867] = 144'hf86fe490f2ba037a14cd1eba0c03154f01c6;
mem[868] = 144'hf4c60fddfa43e81b11811c05e2acec3ce660;
mem[869] = 144'hea9406a41f25eeaa102204fee036ed8d1451;
mem[870] = 144'h03bef14e138519d8e21519eae1fd04fb10aa;
mem[871] = 144'h0437ef0bfe42e0b617d8fa300481efa60880;
mem[872] = 144'he0c4038c009de565f135f492f3e009c2e9e0;
mem[873] = 144'h1296098b0ebae988ec8d1837e9140f0ee1fa;
mem[874] = 144'hfb890847e1c7f21eedeef1dbf5e1ff77020a;
mem[875] = 144'h0c0d0ffaf68508720b8eef53ea9fecdc01e6;
mem[876] = 144'hfaaf1cbf1b20f35006a618b7094f0f931a1d;
mem[877] = 144'h18b403ee1b1411a4ee7afab50455f5d30946;
mem[878] = 144'h16eaf87105201d1cf455e52c04af13b41eee;
mem[879] = 144'he88e0d18e327158108af0df1f94e096eff79;
mem[880] = 144'h061ef46ff4de1f66f717e883078b0606130d;
mem[881] = 144'hed51107801d2fc0df2f4166df0dc1695ebcf;
mem[882] = 144'h1781169608cb1d3be1110033f3a4f0f8f6ba;
mem[883] = 144'h0e0116bafb8305a50f1e101c1a4a00191e5f;
mem[884] = 144'h0b5cf20b0332ed1afa72fd0dea4601b90de4;
mem[885] = 144'h1e0915e61f80f3d9f57b056806a100c60bd5;
mem[886] = 144'hfb46e624065718f80a5cfa3e1ff814691382;
mem[887] = 144'he851f47510bc11031cebea7607ed12080f5a;
mem[888] = 144'hf8b8012819de0f72192e085eee54e870e186;
mem[889] = 144'he0ba0988f79efccb1972ffa8edcdfe19091c;
mem[890] = 144'h05d918fa0a55fbb3fb3fe324e3a80a561b5a;
mem[891] = 144'h0690003ef247ee03eac71236e6d301bde475;
mem[892] = 144'h0ba10069e7a40b2af557ecf80ca413251a4e;
mem[893] = 144'h0a9ff7e1fc4afb56e5a116610b2ff214ec1d;
mem[894] = 144'he33307651f29e40c0281e3f2e23f084509bc;
mem[895] = 144'h00321e51f8331a1e13641c1a16f5f42be4d0;
mem[896] = 144'he4390f22facf1ea7eb311793fdd4f223e02a;
mem[897] = 144'hf6a3f1d6113815acfc141e251d2c16c2f358;
mem[898] = 144'h110a0bf0fd66f1681d62f87cf198f4e6030e;
mem[899] = 144'hfacbe609fe99efc112cb1a39100fe693f245;
mem[900] = 144'h0554f5a60351e32b0d5a17a81571f1f6ef55;
mem[901] = 144'heb5d1a22011cea22fa8fe1d61c49fe10ee23;
mem[902] = 144'h12c903a2ebd6f3721a03120711b606dcf0e5;
mem[903] = 144'h01f9fa2d05afea160184fc3af068130511bb;
mem[904] = 144'h13c7035b0cc7f5631de50d571c131205e52e;
mem[905] = 144'h08a3e8ad0ad4f2cb1eba069b113309cc0420;
mem[906] = 144'h1e2317f3ff61f66ae7b5e490ec8a13c9ef7c;
mem[907] = 144'he076e3f105daec4d12fd04051f80e09bf425;
mem[908] = 144'he7c5eae3090218adecd01fa112f3ec5ae82d;
mem[909] = 144'hedd4f7c904bef7f5f95ded77e129ef87f8ce;
mem[910] = 144'h13eaf32c10b815471f081c8cf67b0bebedcf;
mem[911] = 144'h112810670dcd06670073f87d16bcf220fc74;
mem[912] = 144'h1583fdce0c97f9e3edb90146e86cf80ff82a;
mem[913] = 144'hf50b1aa61c730021f159eabc0843033af6ec;
mem[914] = 144'he89c1d4903660175e4d31e70e8d9e5cb0dc2;
mem[915] = 144'he39203261ba0f974f9ec06f014a3f74d1cbc;
mem[916] = 144'hef63f51211790c50f5421b5503cefa23fa6c;
mem[917] = 144'hfd79e8f409bbe22bec0de5a8e58efd6cf3e8;
mem[918] = 144'hfaa414b41b3cf0d0f7f30062f4dc0e4c132c;
mem[919] = 144'hef19e6630f0b04ec11c5fb44eab4e9fd008a;
mem[920] = 144'h11bef2df01ba073ffbc318eb0a52eb5ae96f;
mem[921] = 144'he3ec19c2ec43e046028800421c10ee2ddfef;
mem[922] = 144'h0bae151714ec14c50c1ae5ac055be9180940;
mem[923] = 144'he6c3150dede21581ed211cfff0c7e927ff32;
mem[924] = 144'h00360834e90c1a19ff5bf6df090bfe8ded89;
mem[925] = 144'h069819cae995ee1a1063ed6c1d191d001a30;
mem[926] = 144'hf2c608c5f249fcf6eec60d3f0c881b74edc3;
mem[927] = 144'hfc7010590d80e48ae46b06f509c51ae6e5d0;
mem[928] = 144'hf959f0aae909e2a014f1e969fab1f900e7a7;
mem[929] = 144'h0550e200e5020d29fd1ee3520531fb96f94f;
mem[930] = 144'he4271f0ae2ef1a42f23a1bf4eaa8e2a0ed04;
mem[931] = 144'h05701a97158413a2e85bfd63ee68148706e2;
mem[932] = 144'hf7fee4440f68f2c503450b9eeb02ef5af286;
mem[933] = 144'h0e46039713fd038f1c4c0018ee681c49e2ed;
mem[934] = 144'hedf40b790a260ab4f088f0cbe2b20f9dfb79;
mem[935] = 144'h16ff0e25076b1e87e283f41eef38f86be196;
mem[936] = 144'hf8f5f89707c1fe16181cfbaef9eb031f1e94;
mem[937] = 144'hfa5814b0f0c61bccf0f1f4cd152a1d6d1f95;
mem[938] = 144'hf997126ae3d8001718f107a51b24e6c30562;
mem[939] = 144'h18fff5da13dd10e109a2f7ce14b904bdf7f4;
mem[940] = 144'h10500cd01f56190ff5aa20241c4b11ad0fe5;
mem[941] = 144'h0f5aecb8f87af11e14e218ba14531978f29a;
mem[942] = 144'hfe4b15edefd5e9b0f544eea6e221ed64e792;
mem[943] = 144'h1b640ef40d0ce133f9fb1eb3fda10b89e790;
mem[944] = 144'h11c5f7171a02f467fdfde0580c630f881c81;
mem[945] = 144'hf7f002f4187be20b1c80eb46e809190e1c8b;
mem[946] = 144'h0b0002391333edbcff281915ff9d10970921;
mem[947] = 144'hf31e0168f28ef351ea36e2f0f8bfe7dc11ae;
mem[948] = 144'hed1ae4f01a170fdd1fc6f6dd1c15f6e2e9b4;
mem[949] = 144'hff70f84dee420ac5e83f1a7d1afb05cdea68;
mem[950] = 144'h0980f0500c7af39e17f7f845fd91079918cf;
mem[951] = 144'h1abd14f2f1ffe069e8971c36e5bff765063d;
mem[952] = 144'h14f6f867e7630fbf16a81da6f9dd07adea9a;
mem[953] = 144'h1bcceee5073de613fcac08e2ef0ef02b1ba9;
mem[954] = 144'he37501a3f589f5d6e9a00b4cf7aa1eb6ef85;
mem[955] = 144'hf1ffeb70e3e1f321f945e367ef75e261045b;
mem[956] = 144'hf1171ddbefbce0c2169dea2317e80fabecda;
mem[957] = 144'h1d21f1750b4b04f71b7ceb13e9521d28112b;
mem[958] = 144'he6851ac71e4d0d76e411e54d0f08faf2ea84;
mem[959] = 144'hf8a00f920415fb07f3b6fa23e432e3e3184f;
mem[960] = 144'he306f0a013d70ba70169f59d1924fb7e0f47;
mem[961] = 144'h1db0100010e2f9fc138719000b66e56dfb02;
mem[962] = 144'hfedc19fb0afa14ea1e1dfc62e58af4cae001;
mem[963] = 144'hfa36e3531d51ff5614440661facb098fe410;
mem[964] = 144'hf08effabfdae02390ab3134e02b3ea84f3d4;
mem[965] = 144'h03f0f3590ae91f2dfe01efd0ecdaea41f911;
mem[966] = 144'h1b92f17f1377089c0fc0fe3e04aaefe011d2;
mem[967] = 144'h05700d30e7d2fb7ee1d1efc016b51306f59b;
mem[968] = 144'hfec3f2bae8a00818ea8c02fbff550c7c0e8e;
mem[969] = 144'he245e95e0aa6fd86e050e229033b1fa01018;
mem[970] = 144'h08d7e0a6fa35191efc69f38eefd414dcebc0;
mem[971] = 144'h1dacf668e6ffe5c4fea2080314310370f865;
mem[972] = 144'hebf212f5167b0ed4078c0ba20f4ce3970554;
mem[973] = 144'hf5dc09931a821562ff5af1d3eb0b1016f7e4;
mem[974] = 144'h0d26f98be1bf111f135e1557f450fbd8f786;
mem[975] = 144'he178e738ec35177419211d87098e058e1f19;
mem[976] = 144'he3dcf086f15408bf1bf11b59e281194be36b;
mem[977] = 144'h1dd7ff3e10500233100408ea032d076712ee;
mem[978] = 144'hffb5fe81ecd2e8da045c10191b51016600d8;
mem[979] = 144'h0583fc380e461201e1f512031be40f2505d5;
mem[980] = 144'h163af812f9a7f4fd18e504e11523e029088a;
mem[981] = 144'h1059100a0121197f168d09d8f36c1dda1936;
mem[982] = 144'hecd0f1b6f84d03dcf10f0e1101bee945f0f3;
mem[983] = 144'hf5d50faffea5fcc214101fe2184df71d1231;
mem[984] = 144'hef33e08dfaa0f33ee1340be9f5411728ee1f;
mem[985] = 144'h11e0130f02b80cc3f8b0e3dc07ba15f80d92;
mem[986] = 144'he5fbf945f415ff641f6a1b0ae8920e41e31e;
mem[987] = 144'h0da5e8b6e923e54902b4fdcf077c1728f94a;
mem[988] = 144'h1c81fa79122013ea1e5b0eedf9a30d75e7aa;
mem[989] = 144'h130a0135eadefdcee5e9f7d1fbe0fdd0e747;
mem[990] = 144'heddbf905fca11e0d027fefabf238ebdfe035;
mem[991] = 144'h081ae7ce116e09c1f973f1f60414ec800c50;
mem[992] = 144'he7d7e37a19ec084d0c670d251f8a000605d1;
mem[993] = 144'hfafaf9730bbff1b0f9e8eb9f01d2f716fcac;
mem[994] = 144'hf41018eee0ecfbeef1711a31e97e1ce70473;
mem[995] = 144'hf4330c3a1754fccc02d0145be6c10d7a198b;
mem[996] = 144'hfb55faa91c691af2f6ee0b89f451fa07e172;
mem[997] = 144'h1def1e59ef06e85eef91e45b0b6f069c0a51;
mem[998] = 144'h12cb0e6cef7de65ef74b0516f054ff11ed28;
mem[999] = 144'h1f9f0f21ffb8e40ff4c4e39e0c36039c18af;
mem[1000] = 144'h116aeecb0d0e1b27f9b600aa1d6e0332f002;
mem[1001] = 144'h0c8619fef912f938033e19441d8a0562009e;
mem[1002] = 144'hf458185803a91d8403bae0c01888eb82017b;
mem[1003] = 144'h1159e3300a9a09c60a1d0fc3f3d80c43e23d;
mem[1004] = 144'h14731113187bed56f81f0588f81ee29ef5c8;
mem[1005] = 144'hec4c17df19fbf558f1f5ea79e4c6dffeeaa6;
mem[1006] = 144'he718e6df0bee1e56ee0ee640e5600f1b1455;
mem[1007] = 144'h080af5acfc0512bc0cd4eb63e98ee45f1117;
mem[1008] = 144'hec9f09020508e6790545f23e1dd01a0c12de;
mem[1009] = 144'hf857e372e660ed6a16f309b50d210cfaf640;
mem[1010] = 144'hf4b4e18710d81805e843f7e4ea450ad1e073;
mem[1011] = 144'he96ef0ba017d155414b4ee470201e6be00a0;
mem[1012] = 144'h0a0c07a9e61f1506fbc70546eee5f1e507f2;
mem[1013] = 144'hf909f6b6fc0ee5a9fb8fe100edc51184f4ed;
mem[1014] = 144'hf9021000f506f8691191fded13d2f8a0f810;
mem[1015] = 144'h0b97e0c4ee8bff4d1a3a1745ef21f9fefb42;
mem[1016] = 144'hfaedebd10d7aff5af5f2e3e2181f1ae6ffdc;
mem[1017] = 144'he0040b201a8818e61911f8c21d2e11ace23b;
mem[1018] = 144'h06d2e121fd170d950175eb44fedde4930a17;
mem[1019] = 144'hff4400a3e764fd51ec7519ade14c1efd1704;
mem[1020] = 144'hf588f7a215e5e9b71411ee18f458ec50e936;
mem[1021] = 144'h0595ff9408190f75e19dea73198cf41af264;
mem[1022] = 144'he112fdcefc7de0701ddbec17ecddf0a9fd51;
mem[1023] = 144'h1be0052ef0f90960e350eaee1ca70311032f;
mem[1024] = 144'hf47118e3ecb7ed721f48e6a10cfae051e7a2;
mem[1025] = 144'h080df473e228fee303f7efceee8b0af21c99;
mem[1026] = 144'h1a31e841045c0d22e9f5e7770df1fe4c1927;
mem[1027] = 144'h1f771959e3630b501cb30ee907c41d5f021c;
mem[1028] = 144'h02000a7703c301790eea1a2e0ceeeb59ecd0;
mem[1029] = 144'h09b9006e0818f70c1fc8013cfd4f056e14e7;
mem[1030] = 144'h0020f6921ee10457166af08f1053e316132f;
mem[1031] = 144'heb790579054be5c21b3e058607701e142033;
mem[1032] = 144'he1ca108f0737e7341021f490004ae457e06f;
mem[1033] = 144'hff33f645f1780758f0c5e86fecf9f1eb1097;
mem[1034] = 144'hf9abe735105b189411f01348f5d1e57cf552;
mem[1035] = 144'h1e8d1314e4d11283f3fc15c30865f6eae58e;
mem[1036] = 144'h17fa1dc5ecc81d5de88ef21bed3d003eec07;
mem[1037] = 144'h194e086dfa4b01c1e38c033fee8fe9b4f292;
mem[1038] = 144'heef306ce0c421015ebae0f45f8ae1a0dec6c;
mem[1039] = 144'he49a077ef6c50c88e52bf1d30e85f6361268;
mem[1040] = 144'h0e7410e30aea10a8130af57e0a27efa2e99f;
mem[1041] = 144'hecb71a8cf148f0200bec06a516491fc5eb89;
mem[1042] = 144'hfcd00f6309deffb0f13401970b2f098c1551;
mem[1043] = 144'he6e0fd6a1d6ee589fd740b5cf1effb1b1319;
mem[1044] = 144'h1bf808acf450e7da1fa6197f0144057bf969;
mem[1045] = 144'he35012ca0a1f16271b3609da01130c3bef42;
mem[1046] = 144'h1a6d1cf3ef77e3330ac3092d0d52e21aef92;
mem[1047] = 144'hef150ca4f0d30e891c45058ff3e60c9214f7;
mem[1048] = 144'hf74e12da1096143ce828f5c1e6d71d8de29b;
mem[1049] = 144'hefb217f4e5a11e690e0d12c7f2b7efceeef4;
mem[1050] = 144'h1bd1ec430c23058418ae168df4ac1285ea8c;
mem[1051] = 144'hed91efa1e7ff0f17ed47f5471eb8fc2506ab;
mem[1052] = 144'h0f3d029c1c09135ce9ebfdd21032e6e3e422;
mem[1053] = 144'h1b46fc62e9defe83f76be0110b611ee01bea;
mem[1054] = 144'hffbffe84e97eec3b107605dbfa2afb1e12e1;
mem[1055] = 144'hfa8ae91517cfe532e7c1e681f58d02e4e511;
mem[1056] = 144'h0353188f158700f8163c04f5059f1072f101;
mem[1057] = 144'h13d9054d042709fc1965fbb5001eecfe0d02;
mem[1058] = 144'h0feaf90708a20707fbc5f5d7f6f20a9b11a0;
mem[1059] = 144'hf565eeda0b061ec5e4731e37eca903d909ed;
mem[1060] = 144'hf557f5c61c77e5e9fe81fd35f2500e2dfdd0;
mem[1061] = 144'h19250bef09b60d10e268f927fb3e14e41a16;
mem[1062] = 144'hf9ef1ce7f93afeb8f1b5e273148c087a11d8;
mem[1063] = 144'h0f23e074e354f513fd03f934fce6105b0838;
mem[1064] = 144'hfbb7f3fa056219c41d790474045817600561;
mem[1065] = 144'h066c047fea510412e35d13d004b5e4d6fef2;
mem[1066] = 144'h1da009130df0fa8ee6ee14020da3f3b4ea97;
mem[1067] = 144'h1f8ae1e2ff1aefaae2f0f314092d1152e659;
mem[1068] = 144'he90df6a9ed31ed86108008ff1cd201b8f2a7;
mem[1069] = 144'h06f515071c42ff25e0a7eaaf151918d000b8;
mem[1070] = 144'h0d121913f3faf49f18e00fa3e0d5ecc9f5af;
mem[1071] = 144'h1496fe0bec750f1e1f3def38e7b9e91fed76;
mem[1072] = 144'hfbdd1c9aeef2f33f060b11591f2cfa3d1091;
mem[1073] = 144'h0f9afe4219890ed3193e089f06f6ff191267;
mem[1074] = 144'hebdbf9310effe4fbf956165de5caeebb1271;
mem[1075] = 144'he26eec8ae4310440016ffa58fa23e652fda3;
mem[1076] = 144'hf7190faa079c0b12f538eba9e1c50e291318;
mem[1077] = 144'h18daf0cc1adcea6f030ef85cff65ee05f2a8;
mem[1078] = 144'h08f00665e1b2e17eedbfe3e2f551f3cef1d8;
mem[1079] = 144'h038d0160f1fafd3bec59ff12ea76e92c126b;
mem[1080] = 144'hff72f8e1f9140878ed03ee32f864e3181848;
mem[1081] = 144'h08c2edcbe21deb60118cef4e004b0877f08c;
mem[1082] = 144'hff0cfe90fee9088308b31503f8f80a71e2ef;
mem[1083] = 144'h10a9e1e6eca01790132fee831415fb70f6b1;
mem[1084] = 144'hede110a8ff8c0ff1074df4aefb00f0e40852;
mem[1085] = 144'h0737f6260e6cecbae76003d311a0167d1eeb;
mem[1086] = 144'hf088f9c2e80d0595faa008b11a9ef83fe634;
mem[1087] = 144'he936f72a16caf97afb60e247f594e656ef68;
mem[1088] = 144'hf40ff2f809cc0c2d0b6f020214c1e5711006;
mem[1089] = 144'hf07ef45ae66de818088fec2603dee43c15d5;
mem[1090] = 144'hf7bbe39de24b10ce14c5eb33fe830a2c0f83;
mem[1091] = 144'he0970389fd43e57df11802911410e5231a05;
mem[1092] = 144'h043f050beb200440e4af09b6f9fdfac8ed0c;
mem[1093] = 144'he589e75cf2f51904f2170682feab10fde376;
mem[1094] = 144'h15b0ea8bf1e100d80c911e0bf5e7164418b2;
mem[1095] = 144'h0cf9f094056dfa4d035af591eb7715f5fc65;
mem[1096] = 144'h1cbd1515e4a31319fec607ef0ac2fd990366;
mem[1097] = 144'h1b12fa8606e7f0f0e5380f49fea0068be2d8;
mem[1098] = 144'he65ff92c1ec4f206f1ac0e99fcc80ff1fa95;
mem[1099] = 144'heb90f3d8f4f715710388f8cb02de0ba8f903;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule