`timescale 1ns/1ns

module wt_mem2 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h08e1f09e05700e080a8707e004070d060739;
mem[1] = 144'hf24208cb021ff1820dbafef800c2f3ecf056;
mem[2] = 144'hf79af41f025bfccd0e04f1d2f2e70e56f74d;
mem[3] = 144'hf6e6f9fef280f3acfd59f82ef95600080970;
mem[4] = 144'h09b6f46b0ef609c304d1046906c7004a0929;
mem[5] = 144'hfc1ff91e0a42028a03b20f71f809f874075e;
mem[6] = 144'h0c7dfd2efa3bef7dfe770909fe4f0835fee4;
mem[7] = 144'hfb780879f5e908340d9df43503db0ee9060c;
mem[8] = 144'h0579ff7b0ab4ffa1f48201b9f5dbf1970d7a;
mem[9] = 144'h01dcf65bf325044f0e1ff450fd2df27ff540;
mem[10] = 144'hf42df22afdf5f6caf7b7f0660ca0f1b80cc2;
mem[11] = 144'h07ad0f0efbb7f7820bbdfbcf0784f2c005db;
mem[12] = 144'hf556f9e80c3ff634f6d20642fa1ff8000199;
mem[13] = 144'h065e013f09cbf4b2058507b80e48f0eff39c;
mem[14] = 144'h06e4fc1e0cd5fad503fc098504a1f06807aa;
mem[15] = 144'hf9cc05f80d47071cf016087308fd0ae7f154;
mem[16] = 144'hffeefa7f0e42063f0a56f09a0ef8073afb6a;
mem[17] = 144'hf6090bdc0d4b06d8026a0961070bf239f919;
mem[18] = 144'h0b7302a0feaa0c83f4adf73d01590cba0cfa;
mem[19] = 144'hf213fdba03650c4e0a570a05f1f1fc840c36;
mem[20] = 144'hf35901e00b5a004cf00f0d75f42308530f84;
mem[21] = 144'hf218f0b40eaefdd70e5d0838f571fda8f006;
mem[22] = 144'h068701240d12f81ff8b0fc4ff01a0de9f055;
mem[23] = 144'hf2dff1e800d2fa4407350a8c005c01cc0b78;
mem[24] = 144'h08f0ff1af236fcbc090602fe069bfb010d80;
mem[25] = 144'hfaad06730e8302fdfc10015a0ca3076c0145;
mem[26] = 144'h0aa90ea00540f178f9070c8c0684f46d0309;
mem[27] = 144'h07f000b403170f26f16b0b36f75c08010f6a;
mem[28] = 144'h08b6f974f8e4fa020220fc3cf68209b00acb;
mem[29] = 144'h0c4a0f9c0cb8f645fcc20fc2fca5051104c2;
mem[30] = 144'hfe35fbdb0a54f5fc0e4703dc08b6f0b40102;
mem[31] = 144'hf4a90a48ff9202b6070404b9f2570d8c0c41;
mem[32] = 144'h0d650ebd0f3e080ef916f971fd7801a9f8a5;
mem[33] = 144'hf26e077f0a08003c00a1f5d5fbbb09b7f3c4;
mem[34] = 144'hf6c207b505c9008bf257f472fdaa0b1e0b92;
mem[35] = 144'h0bf407bafec2fed7fecaffbffdd90b81ff6a;
mem[36] = 144'h04bd07e2f888fecf01a70cb30e04f8d4fe70;
mem[37] = 144'h0b140a6f0d7bfd0e0fb50787fec800c4020b;
mem[38] = 144'h05aef14a098d0733fa11ff360caaefdcfb37;
mem[39] = 144'h0ffd014a0bb80b6f0fb1f203f0f2001e0f5d;
mem[40] = 144'h0b20fb80f800f8b30f30099c0552f28bf2c2;
mem[41] = 144'hfa120948f188070df659097200470579057f;
mem[42] = 144'h05a9fe6df111fbc6f1500e49f25f076c0779;
mem[43] = 144'h0c38f91e0737f08af7eaf66c0ae9ff7df6bb;
mem[44] = 144'h04880d9c0eccf5a702d80c0001fb0a09f699;
mem[45] = 144'hf183f524fa75fbc60cf4f6640897f9fe0870;
mem[46] = 144'hf6b5094b04c4fbe30e7a0c21f7ec038f048b;
mem[47] = 144'hfe070b4600d7000f057a0e8c00c8099bf215;
mem[48] = 144'h052d06d0f747f136ff1304d900c202e7fc1b;
mem[49] = 144'hf91c001cfc2d097f03890750f47a067c0c61;
mem[50] = 144'h0c1d03aa0535f7e5f50001870ec30a32f823;
mem[51] = 144'h059bfba9ffb60339f57afb3efaee094d08b5;
mem[52] = 144'hfc680319fb05f3550f0df81ffd67f6bbf934;
mem[53] = 144'h005a0be7f0a70caaf27809c7f6bffeaef592;
mem[54] = 144'hf33ef18d0b18f5a0f2420fb507cfff95efdb;
mem[55] = 144'hf358f447f03ff6ba0c1cfc0109d70d8af55b;
mem[56] = 144'h042501f0f8f302c9fd640186ffd6f23203fa;
mem[57] = 144'h0a99fc9cfaef080afb62016f03c0f29efe80;
mem[58] = 144'h0c34046cf3b6f17407e9fb3bf2c70ee404fb;
mem[59] = 144'hfe1c0a210ed3f7ac0b090aaf097bfeb7f249;
mem[60] = 144'h06d800ffff2b05bc0ba1fd3cfa12f19f0ce3;
mem[61] = 144'hf3dff88e05b102770181f1bffa7cf5c0f111;
mem[62] = 144'hfb4c0a44f7d5f0bcf82d0513000af17afa92;
mem[63] = 144'h0a04fa95fafa02d8fd03febb00fe093afb97;
mem[64] = 144'hf9430f31074ffbf6fe1800e5f3a0f2e3fb33;
mem[65] = 144'hf0e40f05fc12fdc000b30c3df1300d1bf829;
mem[66] = 144'hf5d4f5f100a6fc5205e60c84fbb102410dcb;
mem[67] = 144'h02aefcc8f818095504f8f100f557f4e10310;
mem[68] = 144'h0167fdaaf83af5e60dd10d230c8cf4aaf8ef;
mem[69] = 144'h0d6600890580f24c06f0fdf00680ffdd0fc2;
mem[70] = 144'h01f1fee6fda3fe8cf2510a03f97ff354f759;
mem[71] = 144'h09f80df20fa903b5f0660449f194f9e202f0;
mem[72] = 144'h0072f8c609e3f2a6f1c1f4440dadf2e9f3e3;
mem[73] = 144'hf9c9fd8201ea07900996026ffa63099af2bd;
mem[74] = 144'hf4b407c4f616015501e20b7e0f6afe670f31;
mem[75] = 144'h01480102f56a0e3f0385f7c202b5fd70fd06;
mem[76] = 144'hfc19f59b0d08048dfe4ef507f3d40702fd3a;
mem[77] = 144'h0f0002700403f11a0412fe5cfff402c307ab;
mem[78] = 144'h09b8f3ec0476f18bf6bb0b24f5bcf3d3f9be;
mem[79] = 144'h0338038af1f7ff5d0e75f785f459055d01ba;
mem[80] = 144'hff660043fca90f7bf9b5fde6f1a1f70d0677;
mem[81] = 144'h0ddbf83bf47d0031f14b0654f0defcb4024d;
mem[82] = 144'hf218f953f7370bf301bf02c102b9fd81fcca;
mem[83] = 144'hf9fefbeff53500c8024d0da8fd9b0ec70e5d;
mem[84] = 144'h0819f8db0e71f67202e70e6b02ddff100d2e;
mem[85] = 144'hff71066d073501b00cd70b66f7300b78f5cc;
mem[86] = 144'h0961040df9b2f96cfb2dfd570604fe8bf083;
mem[87] = 144'h0eac0e0ffdf8f331f9e80d270f14039ef58a;
mem[88] = 144'h068c00ab0ee50fc50c1c00960c5908ad0bde;
mem[89] = 144'hfa680f96fb44fca5f3e60051f1290f85fd73;
mem[90] = 144'hfa42fda8f668f712f3de0c8502d0f75bfb6b;
mem[91] = 144'hf273f056036bf26dfa17f2f4fc99f7f60d87;
mem[92] = 144'h0d8f0bbbfccff139f8cffdf20b1f081bf812;
mem[93] = 144'hf3070a68f9ae01010d460f0c042c081501f4;
mem[94] = 144'hf5d5f0a3028cfef5f0910756062b0a5e0007;
mem[95] = 144'hf20707b5f402020808c80e7af5cb05c50459;
mem[96] = 144'h0cc6027308d40383f9140433f0ac0a9bfc52;
mem[97] = 144'h0413f88af70e0d9703c6090b062c06dcf923;
mem[98] = 144'h037bfec3020ff99cf0310e09f5da06e8fc11;
mem[99] = 144'h0579fe2d0403031afcb1f162fa750beafcea;
mem[100] = 144'h0c120f4cf171f439003300850a160750f1c8;
mem[101] = 144'hf22d08dff6edfd50f610f7a70fac02edfebc;
mem[102] = 144'hf08cf6a302c80ad0fb2106fc03cff66dfe9d;
mem[103] = 144'h0815fd24f4d7fcc60edf039af0280658f686;
mem[104] = 144'hf147098c0a57fde9ffb5ff73069bfda60958;
mem[105] = 144'h0dfdfde5f180f6dd07d00455003e068af1be;
mem[106] = 144'hff51f942ff5f0e36f8400824fa6bff0c0bb0;
mem[107] = 144'h0e170ca40d80022703070d47fa890c78f7d7;
mem[108] = 144'h02b605c9048df3ddf7e5f646f2070537ff84;
mem[109] = 144'hf6defa8effbbff5cf0270a710f3f0069f387;
mem[110] = 144'hfee8f62b0893f823f94afa83f9720f54068f;
mem[111] = 144'h02d402640fbaf8bd06e80977f1f1f2a9fcd2;
mem[112] = 144'h06660890f04b072109790a5f058f08620bdd;
mem[113] = 144'h01960b06fdc6f0150589095ff80002ab0a18;
mem[114] = 144'h0660fade0fe1fccdf93503c4f26ff25602f8;
mem[115] = 144'hfc9dfbfaf806f6cf0dbbff3a0226ffa1f150;
mem[116] = 144'h0c990eacf0730a4ff6fd06a001c1fc75038d;
mem[117] = 144'hfaf8f82dfc42f6fe0cae0afcf33c047501d0;
mem[118] = 144'h0772fca0f851facdf3e10abef33ff9110634;
mem[119] = 144'hffb4f9610c550f130b250e1f0053f9330c82;
mem[120] = 144'hf74b0fb80c43f825fafbfeaffdf6fc5a0b4f;
mem[121] = 144'h0bc40930f06af507ff5f0a1809b8fbdd0fd9;
mem[122] = 144'h0906f85df77ffedd0b2f095c0fc5f8aef29c;
mem[123] = 144'hf04bf2240998fefc00cdf3c9058ef6bcf162;
mem[124] = 144'hfb1b09870a01f9670b310b810b55026a0c92;
mem[125] = 144'hf2c1f08107b7ff7af434f66608c201c20508;
mem[126] = 144'h005ff97ff51b0ee5081ef291fe1c06ce09f6;
mem[127] = 144'hfc900076082f0baa0ce8fca70285039a0ef6;
mem[128] = 144'hf3a70e1bfe94099c0c7af66bfa26f012f0b9;
mem[129] = 144'h0659f0d0f5f1f14bf537f4fff1490ddff0cf;
mem[130] = 144'hf392fa2ef438006afc03f805f4e802ddf1f9;
mem[131] = 144'hf705f253f861fba7fb90fc2f0a76fcf1f949;
mem[132] = 144'h0b62074cf2d107870e77098f0a10f4fc020b;
mem[133] = 144'h01480d43fb0eff490a57fbca0a2df1d10503;
mem[134] = 144'hfcd8f59407a90f8dffe70539f928fb0b06ca;
mem[135] = 144'h02eff005f53304aaf307f82cf4a5f5f60c19;
mem[136] = 144'h0a8e05a6025807550a3a07a90a0e0d6f0a81;
mem[137] = 144'h043801750dc1031c0ff209240df10687f619;
mem[138] = 144'h0eb00fbbf570fec8f5aef446fd7bfb250beb;
mem[139] = 144'h045df9b4fa2ff1eafe3ef53305a803de0f35;
mem[140] = 144'hf97c08c3008905b802e0f8e1f1d4078d0498;
mem[141] = 144'hf284058107ebf07206f6fbd9f267f92705a6;
mem[142] = 144'h0db006d1f8cf0813fc2d07acfcba06d4090d;
mem[143] = 144'h0efe027cf061031d024ef60af21df4a2feea;
mem[144] = 144'hf9e1f9e20152f17a050cfd1406740e0bf088;
mem[145] = 144'hf80000d3ff0c0939037e0a1bf975059ffdb4;
mem[146] = 144'hf310feb70e8cf1faf4b0f3470a750b95f691;
mem[147] = 144'hf7b4fe100adaf9830e520110fc88f40cf105;
mem[148] = 144'h05dd073100920c97fb97f663f13af4870562;
mem[149] = 144'h035cfa790ae8fffa053bf08405e7ff7609ea;
mem[150] = 144'h06ae025bf712fce1fdd501a8033b0365fea9;
mem[151] = 144'hfbe9fb38f00e090df153f647011d00cbf5e9;
mem[152] = 144'hfef0f6430d6afc5b0e3effd30b4700c80f57;
mem[153] = 144'h01cb0b82fe27f467fedcfd4cff6809a0f87b;
mem[154] = 144'hff46fa130de0f26a0e46f8c9f867fba30832;
mem[155] = 144'h0dcd0cfff83cf378f3c80b22fbc8fbac0c04;
mem[156] = 144'hfadbfdb3f045049401b706350f7008210eb9;
mem[157] = 144'h01cff775f9fef23c09b7fdb806c108c9f73c;
mem[158] = 144'h019d008af21ef21ffbd006b80c5df764f58a;
mem[159] = 144'h019501370c3e041ffd280723fc4a0d3ef75d;
mem[160] = 144'h05ee024d02d704f403760eb8f018f4abfa8d;
mem[161] = 144'hfb6ff62e002c02980a4b07a8f2e90db30c7a;
mem[162] = 144'h0321f78cf3f6f767f260017af9a1fe540717;
mem[163] = 144'hfc5d034dfc8a0b38f0ed0fc703e20d890b7a;
mem[164] = 144'hfd0204a30c1ef518feacf36b0b250cf1fabb;
mem[165] = 144'h08d2f5770efa032e04f407a7fc82f3f408ab;
mem[166] = 144'h0464f89eefc80097f73a0e7a0bb004c7f2e3;
mem[167] = 144'hf486ffd70b85f2650ce0fe120c6ef8aff97d;
mem[168] = 144'hfbd2f439f2e902a80492f4c9f5c0f6c3fa34;
mem[169] = 144'hfba30cc00638f0290129f8b4fed0f29ff34e;
mem[170] = 144'h0034f80905bdf92d0c060df90b7104fcfccb;
mem[171] = 144'h0026f11ff821f2640b2105bcfe4e0db20922;
mem[172] = 144'h0439f16e0feef5d9f673fabefff8f8890590;
mem[173] = 144'hf2bb0b8206f802040a310cf9f090fdf30280;
mem[174] = 144'h0069ff9bf27efd91f02cfdd0fb61064e0549;
mem[175] = 144'hff29f55a0552f4da0188f0ad05f1098af3b8;
mem[176] = 144'hffeef34cff8cf499f0fbf20b0e9f0b4e05ac;
mem[177] = 144'hfe61f94a0f75fcfbf93902aa061ef63bff06;
mem[178] = 144'h09ecf0a7f5bbf3c9feb5fe01fc3904d50267;
mem[179] = 144'hf0fdf98cf3560f23fde10cd60eddf02cfdd7;
mem[180] = 144'hf182f2bffcdcfd830a9503cbf3a5fb45f131;
mem[181] = 144'h04f7f727f901f92000dff5420c65054bf941;
mem[182] = 144'h0485f2ceefd6fffef5e20c9309f60f41048d;
mem[183] = 144'hf93af29c0f25ff4c019d0be7fe72fe2dfaf3;
mem[184] = 144'hfd890219f2c108c30f00056efb30f8f6f79e;
mem[185] = 144'h00de08fa0e0d0a4bf29005090addf1fd0e2e;
mem[186] = 144'h0268fdff08090a7b06360f9f030ff8da03a7;
mem[187] = 144'h089805c9ff0bfba6fd480d8c060508b304c7;
mem[188] = 144'hf4690400099cfd560ac304cbfdfa0d540938;
mem[189] = 144'hfb060b16fcb40e87fa750eb1f7600b400ee3;
mem[190] = 144'hfc500d32078c066ffa66f692f5cef1950c9a;
mem[191] = 144'h01d60c990a06f895f689f0120ef3eff505e5;
mem[192] = 144'h04ef0ad3f8e30036f4fbfd23f2240c7f0ef6;
mem[193] = 144'h09090f7cfdfdf151f6ab031df9310e2bf69d;
mem[194] = 144'h0a11051004b0f329fbd4061e04d2f9b1f662;
mem[195] = 144'hfb18fcfdf62d03da0652f0600a82f5f0f2eb;
mem[196] = 144'hf79f00e201f60420094df0b6f4d4f51af925;
mem[197] = 144'h04f9f46a0f150123f4a6f081fc380873f5a9;
mem[198] = 144'h0ea3f8320d6d0220f80df3d8fbf5fd6b03e3;
mem[199] = 144'h044bf58406f5f1f90ad8fb24f54ef126f589;
mem[200] = 144'h01e5f32b06520699000909c7020af8d1f5e6;
mem[201] = 144'h062e0c1af063f5db0ef00092f3c2089d04e2;
mem[202] = 144'h08380c71ff30031cfd6c0e60f010f1e2058a;
mem[203] = 144'h017bf878fe2f046ff174043cfb0a0089f3f5;
mem[204] = 144'h08e4f20806a508ef0355fe2bfdec091bfcee;
mem[205] = 144'h014d0f2b00d3086efa3e017e070705b6f6d2;
mem[206] = 144'hf60303b3f362020ff2720c210d590488ff75;
mem[207] = 144'hf04108b1fef50dde084efb36fbbf07a8fd77;
mem[208] = 144'h0d0bf1defcf9f276064408ef06fc0d30097e;
mem[209] = 144'h0cd305a106b3fe0a078cf0d3f198fda3fb46;
mem[210] = 144'hf2dbf512f4120c790a5e08490a26036c0af4;
mem[211] = 144'h01a9f32dfb610c80066f08d90a06fa48f445;
mem[212] = 144'hf0630b3c03200314fe1cf13307470be00dc7;
mem[213] = 144'h0251023c0311007f037b0282fe13f3c00ac4;
mem[214] = 144'h00670a7bf0e80c5df2b7fe38ff590a74f47d;
mem[215] = 144'hfe32046506fefdd8f9d4f33afbd20dc6f58f;
mem[216] = 144'hfeee0a54f3e30e310caf044bf5c1f2edf06e;
mem[217] = 144'h0759f2fcf830f26803b1f116f4aa0b7c0be1;
mem[218] = 144'h0909f2710e21f98a03dffffb0b65fbc70b61;
mem[219] = 144'hf745f57a0a37047d0218013ff47609effdef;
mem[220] = 144'hf8e002640482f36208dc075ff94d0e76fb27;
mem[221] = 144'hfa770a04f5590f06f4a3faa30ba700ba074f;
mem[222] = 144'hfdb90439002bf509fe3f0de7f00af5410fc1;
mem[223] = 144'hf9ca07dc0bab0154fb850d460dc8eff1efe5;
mem[224] = 144'hf807f2eb0b8401ef0d67018efe800cd1029f;
mem[225] = 144'h050605db0dfff9be0f8e069ff130f69e0b21;
mem[226] = 144'h076609aff29af1110133fcc80885f8ecfd8f;
mem[227] = 144'h01deff420bfc0f630053ff870e90f19bf7be;
mem[228] = 144'hfc36f6b8f266f97603f8f3b1f67609b80998;
mem[229] = 144'hf932048cf5fbff4dfbf709920bea06fa04f1;
mem[230] = 144'hf0690818012ffbfff8a0f9b508e3f610f677;
mem[231] = 144'h0bbd0dbc0199017900a40878f890f3c70901;
mem[232] = 144'hf64c0a3104460852016dfe18fee6fc0df884;
mem[233] = 144'h0491f739ff43f2e9fe6405ab0544fb510d30;
mem[234] = 144'hf729fa190589f4740e4a042af049f86607c4;
mem[235] = 144'hfbc206beffe20684f3450bbcfba404e3f019;
mem[236] = 144'hf978f53100e7fd3df55e004efa5109fdf9ae;
mem[237] = 144'h03dcf1930644f78ff9220c50f7bcf0c90e3d;
mem[238] = 144'hf7f202bff6b708cafa31f7eb0029fbba0470;
mem[239] = 144'hf81f05dcfaff0f17017b011c0ce20b81024e;
mem[240] = 144'h03c407a2fe77f662011d05e5f771f7a30708;
mem[241] = 144'hfb070bdcf63808030655f4750f78f993f43c;
mem[242] = 144'h0cecfd1305180ad90a290228fbf90996016e;
mem[243] = 144'hf223f95b033104b30385fc7cf5dcf4a0f721;
mem[244] = 144'h0d070a74fc8709060e930a32079d077efa98;
mem[245] = 144'h08dff7cffe9a0273fddb05b30c5205dd0368;
mem[246] = 144'h0a82fb78f5e80ec0f60ff3f5f701fc5904fa;
mem[247] = 144'h06120a8a030d0b3ff63d0ca20f6e009d0578;
mem[248] = 144'h0aee08a40f13f55f0a25f849f5dd073ef857;
mem[249] = 144'h0880049501f307f90cf0f8940a0705c8f0d4;
mem[250] = 144'hf50a0d6aff3dfbe5fe37f09309cbfd750b24;
mem[251] = 144'hfcbffc49012d0fb4f4e5fb6509300d4b043e;
mem[252] = 144'hfca306d7fb6508d6f34c06bc0f9400560a14;
mem[253] = 144'hfe5c0c4bfa78fad6fcf7066ff43d06a0f13b;
mem[254] = 144'hfe300ea0fad7f1a10d53031b0b5d04aa0990;
mem[255] = 144'h0a88f34101c0fa58f3990d79f855fc84f45b;
mem[256] = 144'hf933fd2f07f9fa1c0c880199f3ed0df00ead;
mem[257] = 144'h0f4df7f0f568f072f1cc0d96f18af29406c9;
mem[258] = 144'hfe78fa79f0e0003bfebbf694f613097000dc;
mem[259] = 144'h029ff06bf825097907cc0a2d057407430baa;
mem[260] = 144'hf9aff69afb5cfc36053bfc0f0bbfffbf0796;
mem[261] = 144'h008002aaf3c2fc6202f4f951f689f0ecff2e;
mem[262] = 144'h03df02f0f501fb15fd21fa05f4dc01c4fa50;
mem[263] = 144'h0318faa4f32afc53f032f5d00c8c08d40113;
mem[264] = 144'h020f084df9ebffcd0bb0029202ccfd050d1f;
mem[265] = 144'hf6f7fee008150d660cc7fb7409ce0321fe6f;
mem[266] = 144'h02bff8ccf59dfc120f9ffbe8f068f65bff8f;
mem[267] = 144'h086afc76f5f4f22b00a105e70e1c0c3404a6;
mem[268] = 144'hfa15fbfc06b9fde40101fed80fdd06fe0082;
mem[269] = 144'h06c0fad209e60b240df30f4c09b50e38fc1c;
mem[270] = 144'h0d67030ffa52eff10172041ff8370758f3d2;
mem[271] = 144'h0a5809f805a1f0b8ff0df637030ff08504e6;
mem[272] = 144'hf75b0c4c032e0b9af20a0b6afb220e44f878;
mem[273] = 144'h01bcf0c804e7071209870d91fe00f7800be3;
mem[274] = 144'hf23d07df0f83f37cf0420e30048f0e4bf5b0;
mem[275] = 144'hff330c42fb3cfcd2099d0bbe0781ff320838;
mem[276] = 144'h0b9eff31f7d50f69f887f755f6aafcd80228;
mem[277] = 144'hff03fb4e06270d3b0c1100d8093b0d860374;
mem[278] = 144'h0343faa405a5f5b7f02efb50f7aa0e4cf88d;
mem[279] = 144'hfc49f0a205ce0a4e0e10058703f2fa2e03b3;
mem[280] = 144'hfbc207dd01f5f9390a0af9b908c4f76cff38;
mem[281] = 144'hfd970638f7cbf35bf3e409920baff605fd62;
mem[282] = 144'h008503f005450e6e0aa3f04a015608c8f2b9;
mem[283] = 144'hf669014c0461feb608d60509f25ffd26f532;
mem[284] = 144'hf741f6ee0e6ffc320a84fe37f21c0807f651;
mem[285] = 144'h02d7f26afa3cf1fb00b10e26056df7670782;
mem[286] = 144'hfb0f0883f4d80c3bf954f155ff64f0e30dc7;
mem[287] = 144'hf0b6043208fbf502f4b1f6580262f7caf51b;
mem[288] = 144'hfa46f414fa45f52ffd92fa1b060d0f09f315;
mem[289] = 144'hfabb0c750688f45a0996f9790204f95ff3ae;
mem[290] = 144'hf7b807e20142ffb1f0280067f01dfe30f288;
mem[291] = 144'h052ef6a80c43ff67fac60fd80a39fac4faec;
mem[292] = 144'hf4a9f999f374f6870724fbc707510b9af083;
mem[293] = 144'hf3f40704081f05a4f3b5f572061800f1fc18;
mem[294] = 144'h0685fdd5053d0213f6100b390f35f14dfd0e;
mem[295] = 144'hff15f7440a69f83f01030082f9da03baf864;
mem[296] = 144'hf2f7f802f9a70b9808dd0a3b04e401a70fe2;
mem[297] = 144'hf8f8f4bbfcd3041ef8380e4bfd0e04adff8d;
mem[298] = 144'h0b20ffb2fd4b0c1cff82017efcb5f442fd7e;
mem[299] = 144'hf833ffac01d8f14007d2f5290cb20bab0d71;
mem[300] = 144'hf77b0e1c0901f18101240160fd6e044cfcd1;
mem[301] = 144'h04d40d7dfb5201c4fa5809f90868f36a0dfc;
mem[302] = 144'h0fbbf9a1f634f287f16e02a2017f0e16fc35;
mem[303] = 144'hfb90075f0028fd590c6ef5740ba3038b0762;
mem[304] = 144'h010bf97bfc29090ff9fef6b4f4980f83f59e;
mem[305] = 144'h03c1fcc9f0dd096dfced0166039700da0ed6;
mem[306] = 144'h076bf558fbcc032df551f8b2f90dfe9efed9;
mem[307] = 144'h092705a90cc0f20b01ddf63e05caf793fc50;
mem[308] = 144'hf9e0faf0f39708f301f4f595038df5c1fd9c;
mem[309] = 144'h0adffabdff5bf9510f56010b03d4f6770b84;
mem[310] = 144'h00fbf821093b0640f879f5c90146f1fc0b26;
mem[311] = 144'hf93c048e0937f1a0f3190b6301def262f9fb;
mem[312] = 144'hfc0909fefad9055d0c12fa7ff1c0f1d3f0d0;
mem[313] = 144'h0a65f66df27c0a69032cfc67f3b0fa830ce8;
mem[314] = 144'h01d60003f401f67d0d20fd48f93bfaf3f800;
mem[315] = 144'h0d270281f80205030ced0f02098df354f4f5;
mem[316] = 144'hfbf5f2960ba2f2d807a6f2d90151f547f795;
mem[317] = 144'h0e7b0b6dfce8058e0eabff22f9bcf0faf537;
mem[318] = 144'h08ec0b17fc09fb40f13902e6f41bf52804c5;
mem[319] = 144'hffc5f1220ab1f9e2004bfb98fe03f43a02a3;
mem[320] = 144'h05fc0bca0f9107700131fcc509490a38fbeb;
mem[321] = 144'hf629fa050bb6055009d9f6bbfaf3f36df419;
mem[322] = 144'hf14af3c00683f2e0fbb1f752046f0330f0f7;
mem[323] = 144'hf612f4e9fe1d09900b240b9cfa8ffe6b0306;
mem[324] = 144'hfd5b0da6f88b0b0a0f2208ca00680d98f0ec;
mem[325] = 144'hf4bfff0f059f0e980b2cf68bfcb70203ff21;
mem[326] = 144'hf1ddfd8c00420022029df2ec051a0cd0f96e;
mem[327] = 144'h0ef3012ef2fb0d04fe35f94e088af1040b12;
mem[328] = 144'hf233fd5f03dd05acf0bb01a605f5f3280c24;
mem[329] = 144'h01eefbd1f638f295f5c30efdf098fd530ca4;
mem[330] = 144'hf832fa8605c8f2c2f65a08ea009dfa070371;
mem[331] = 144'h051bff18f6d1063bf6d9ff430778f02a026f;
mem[332] = 144'hf244f3710fe6f2c9f476f04df9b1f914fc9a;
mem[333] = 144'hfac40a030f11ff6a0a0c02c500d7f3dffad9;
mem[334] = 144'h0bf1f070f2cf08aa079dfc02f826f079f66f;
mem[335] = 144'h0f84f16f0981f9d209c7f4a40cfbfe0cf038;
mem[336] = 144'hfc2c046c0934fe2e068c0a0b0831f78f0b97;
mem[337] = 144'h05bd065efa48fed70d5b083d0ceafec9f923;
mem[338] = 144'hfd95f5910e510f4c06fb0e7e02f20af6fdeb;
mem[339] = 144'h0ec40f2df89afb2402c3f9d5f11cf5ef011e;
mem[340] = 144'hf6b9f0f6f882fec2f9a0fa8f0eb20a4e0913;
mem[341] = 144'h0888f72106eef07afdfe05e1f4ac060dfeba;
mem[342] = 144'h01c7f118095b067af397f0880589062d0838;
mem[343] = 144'hf289f8ec0d2f069407f3f9a5f292f24df1c8;
mem[344] = 144'hf6200bc40b8af3970f560cf80527fbfbfef1;
mem[345] = 144'h08d3fa8e0c5ef085f85ff31ff47009d30405;
mem[346] = 144'h00c2f07e01ecfea6ff93089efe700c1f0b76;
mem[347] = 144'h0886f4080832f38dfc9ff7b2f90e067f05b2;
mem[348] = 144'h099e0bf80cf2f59cf4ab02fbf863fc9806f5;
mem[349] = 144'h0e43f872f65204c50e7df74402580ef502a7;
mem[350] = 144'h03140b5902a7f24bfb3d0cb3fab9036df3bc;
mem[351] = 144'hf3550ce60c36f2850e310dd0f67f0933fbd6;
mem[352] = 144'h081708f6fdbe0edafb140475002dfbf6f883;
mem[353] = 144'h07d30a8605f2fc9bfe88045af5c104290a43;
mem[354] = 144'h01490413fc3b04e5f519060ffa68f0fd01d9;
mem[355] = 144'h011f001301b60b2d0043fd26f3d8fa5dfa8d;
mem[356] = 144'h088e070a0df405bbffe7fa1af5e605f80f62;
mem[357] = 144'hf186fd83f6c3f71b0a9cfc6bf17bf876f9a6;
mem[358] = 144'hf21bf27b02810d02f4eb098403a20b43017e;
mem[359] = 144'hfdb2fba5fb8c05d60105f713074a0b37fac3;
mem[360] = 144'h0e46f4a0f71a03830c1af1d7f19c0e71f4f8;
mem[361] = 144'hfce1fb1d050b0cc7f58f0d8605a906b10bb0;
mem[362] = 144'hf825039f0cadf3e50335f4bc0d1101840673;
mem[363] = 144'hf4960a19f03c02adf486ffb0061ef3120cee;
mem[364] = 144'hf7470851012a03ab0da3082ffb37079cfd51;
mem[365] = 144'h07e7087ef332f688fd42fe4b09740084f9d4;
mem[366] = 144'hf33b0b94f687ff70f88c05d203a30003f7fd;
mem[367] = 144'h0e2dfeabf6190f1301ce010dffe70a5f0945;
mem[368] = 144'h0e9201980b01f04bf01cfbf70d040d06025d;
mem[369] = 144'h0ff4fe8dffe1087604f10175f9b70b730afe;
mem[370] = 144'h0e850af0062bfec1f8eb06a60fa5f5fe0470;
mem[371] = 144'h0d430c7ff5ae0fbc0b4e0a1ef914f8720b4c;
mem[372] = 144'hf7c2fc08f5f50982f916072ff66cff030614;
mem[373] = 144'h085e03dcf4610a6af95df756f7d1fdda01a4;
mem[374] = 144'h080cfab700700c07fd7af830f21d08a708c7;
mem[375] = 144'hf29b0314fa6308530db2f479fe7c09df0e1a;
mem[376] = 144'h09b80e54fc25fb9604b805bb0861f2b504d1;
mem[377] = 144'h05ee03920439ff5d0045f01f0aecf99a0552;
mem[378] = 144'hf47f0f72f86b09d001d6f4cff181f1d004d6;
mem[379] = 144'h0090f0f8f4730d69f7550bc6f3190c3e057c;
mem[380] = 144'hf629f2f20ded050a04d4f566085c029103bc;
mem[381] = 144'h0d26f5990630f5e5f43d018e0b5f02d10bbc;
mem[382] = 144'h0da4ff630de8fbc00c2f0af10a20fa78f44a;
mem[383] = 144'hf898fb2cf25b006b098d0096f19afe3efcaf;
mem[384] = 144'h0acdfb62facc02d7f3fafae8fafef109f371;
mem[385] = 144'hf5d80506096df3d6f90a0cd8075507e90918;
mem[386] = 144'hf6af004c03440ba304a204fef3f10e31f118;
mem[387] = 144'h04a9073a0b58ff7b05e2fbad0ad20a8bf846;
mem[388] = 144'h0c4302c8003cf789f25f02b704f50c6908f3;
mem[389] = 144'hfb36f2e8ff3108e700600261f5800901025e;
mem[390] = 144'hf11af68dfc81f8d8f1bdfb5efeb70e7808f9;
mem[391] = 144'h0b4a0aa10e9bf0fafc920eaff4a2fa2af42a;
mem[392] = 144'hf3e4f4e2f6f8fd0a06a6069cf0ef0cd8fb4c;
mem[393] = 144'h0a900032f0710a1204170a2f0356f32dfb3c;
mem[394] = 144'hf0f50335029bf4940bc700f7fb5e09fd091b;
mem[395] = 144'hf762f79cf1420e08fbc90a040f6208db01f0;
mem[396] = 144'hf83102f30c7ff44e0c52f68cf58ef14bf669;
mem[397] = 144'hf6f50139f1610bbbffd203fe0680075701f7;
mem[398] = 144'hf92106750b1708ae07ca0bdafddb0c31f4de;
mem[399] = 144'hfc2ef8670142f6540c4dfc3907230bbefe52;
mem[400] = 144'h0a02fff0f2c8fc71ff01f7260871f66fface;
mem[401] = 144'hf0f0fbb90d20fc7af0da095df264f53a034c;
mem[402] = 144'hf3b4f54808b8f863f92f08e2078b0e5406ad;
mem[403] = 144'hf4e5ffb1f730fb63f349fd670cd7063e0dcf;
mem[404] = 144'hf966fa88f4b00809f39008e307a30f54031b;
mem[405] = 144'hfe80f4b80fe8f9a407c7f3f1f8170d51f46c;
mem[406] = 144'h0e7c076e02380d59fecf0980fb27fbf20def;
mem[407] = 144'h0c1906dcf2e403ccf4e4058ef29606e6080f;
mem[408] = 144'h0eaef115fe14f6140e090e1b0c89ffccf2f2;
mem[409] = 144'h09c6f81ef5df0d9bfcfe0bbbf53dfb03f6f4;
mem[410] = 144'h061800560225f729078901f0f6ac0513fd47;
mem[411] = 144'hfbb1f7e5056efe61f75ff9fa0c9505acf08c;
mem[412] = 144'hf26006970219068100980c70effdf14bf11a;
mem[413] = 144'h04020a91028cf07ffad600c4f1b800a80f11;
mem[414] = 144'hf97f0898f5820a9f0dea001ff05f0edaff30;
mem[415] = 144'h04b0f4550653f72dfcec018108e4f672fb05;
mem[416] = 144'h0bd6fdf605d90e51fc37076f03a2f9e7f1e5;
mem[417] = 144'hf72e0fdd0890f6f10e9b04fef279f0de0340;
mem[418] = 144'h04ad06db02f00a5dfa4d0293f503fe7ef56b;
mem[419] = 144'hf1ab036ef561f1bd0010f2ebfe65faacfc79;
mem[420] = 144'hf61a0bad0d760d71f268fb81fbfaf108f91b;
mem[421] = 144'hf18df4c80c2f0bacfc2bf91d0e9dfc9b0714;
mem[422] = 144'hfbf6fff1ffc6f60f0e6f021e035dfd79f39a;
mem[423] = 144'hf73df43b081f00890b1609c00cb30b24f221;
mem[424] = 144'h034bfc63ffcf0a93fdd30ea106a1f825fb64;
mem[425] = 144'h0afb0fc6f0cbf46cf30108ea022b0ba7f578;
mem[426] = 144'h0252ffcef225069ffa67f9fdf602f3bff399;
mem[427] = 144'h0dec0cb5f8b60f8d02800df60b0ffd7b0850;
mem[428] = 144'h0812ff5801290f34fcfe017dffabf3d001d0;
mem[429] = 144'h0bc1f5f3f696f75cf1ac016ff9080e57f76c;
mem[430] = 144'hfe0af228056e0126fd53f2edf5f0f29bfeed;
mem[431] = 144'hf52c08c8f0770561f33cfebef58cf4830d75;
mem[432] = 144'h057300eaf064f75cf5a7f09d05aa095104f0;
mem[433] = 144'hf392f649f2cc0637082af21e0749fb15f97d;
mem[434] = 144'hf3760d00fc08fa78f4eb001afde509df02eb;
mem[435] = 144'hf075fb22f0d90d29f07305530fa1027d05bd;
mem[436] = 144'h072a0b560db60fd40fe0f5e90f3c0a5e07db;
mem[437] = 144'hf962f2caf10a0d9bf84ef24b037afc6cf650;
mem[438] = 144'h0fd1f21101b0f76a0c4808e5037df8260b88;
mem[439] = 144'hff2ef6fffbdc0210f5340107fe62f1d40e37;
mem[440] = 144'h0596f92008450e0d0cfe0a04f2baf96b0512;
mem[441] = 144'hfb0300e60937f479faf90cd10ae30c0aeff6;
mem[442] = 144'h00e8f6a2058708cef152f68bf692f8cd0975;
mem[443] = 144'h0310ffce047d0ac800d5046c04a70e65fc75;
mem[444] = 144'hf7050cee00cdf4d30a6f09cdf8dc0c14f198;
mem[445] = 144'h0df20f7300ad08a3083d0116fab9fc0e0b31;
mem[446] = 144'h0c66f5980e25f153f2ec083f0582f06c0762;
mem[447] = 144'hf36109c1fe640477fb06f185076df37906a5;
mem[448] = 144'hf2e604cc04a1fdf30a4af38e01e3fa720235;
mem[449] = 144'h02b904a5fa69f7b303a1ff65f75909e20d8b;
mem[450] = 144'h0f74f6fb0b380e1ffc670c1d0aa00db80374;
mem[451] = 144'hf64400cdfa4a0666fe04074bf114f931f8c5;
mem[452] = 144'h0e9d0187f45f0c41032f025bf12005190634;
mem[453] = 144'h07d905990e2907cff82efc39036a0519f8ba;
mem[454] = 144'h082dfc4c0b1c00fb0cebff60f9a1ffbd0af3;
mem[455] = 144'h0438f6b5f29b02570b1d0a170c3504fe04ae;
mem[456] = 144'hf7acfaa4f4ac0ca40f3a0b70fa8e0326f486;
mem[457] = 144'h0dd0f9c9f9690bb900b2fb0bfc2c0f24ff67;
mem[458] = 144'hf62b045ff02705ecfb5303d0f3ad00f3faf9;
mem[459] = 144'hf4eefb0ef541fc39fa71002f05b2ff5ffe21;
mem[460] = 144'h03c9f2c7069cf2f4f942feedfd49f731fdc2;
mem[461] = 144'hfce60a8607e5fe22ff7bf848f69d01e0fd08;
mem[462] = 144'h0246ff64f26ff7e4fcb401f705e20d51028e;
mem[463] = 144'h0e25f648f7990fc00788fa13f978035502f9;
mem[464] = 144'hf0dd0da9fb560d540a45f848f8380619ff83;
mem[465] = 144'hf812f1a0fdfc09920c8cf799fcba0ecd0b11;
mem[466] = 144'hf7f20bc6f736f7cf0ca4fc82fb84058408b7;
mem[467] = 144'h00e30970019bfdde0ce2f9810b80f870f0c9;
mem[468] = 144'h0cc2f1520be3001b093fff75fa70fe58fe29;
mem[469] = 144'h0d9401a10c63fe02028b0bc7f8000e630624;
mem[470] = 144'hf298f81105dcf421f6d5fdf50ad2f032f922;
mem[471] = 144'hfceef8160f44f6ab0adbf84dfce00a26f335;
mem[472] = 144'h0dc904e10c49032cfdeff54ef454f4610727;
mem[473] = 144'hf244fceaff6cf9c40fb60bba0387fdbaff30;
mem[474] = 144'hfe7f0778025ff3c5081ffea8fb2407650679;
mem[475] = 144'hfe5e0d48f8ae0c16f755f463fea20903f72d;
mem[476] = 144'hf285f960f033f744f532f16f0c520c86fd90;
mem[477] = 144'hf1b8012dfc5700aef549f533085df317fb44;
mem[478] = 144'hf9a30b410281f42cf3650068f49ef869fa6d;
mem[479] = 144'h094a0c570b6703e1fd79fb1efa0bfb5a0b9f;
mem[480] = 144'h09a3efe2fa4e089af4eb03760eb4fe8ff6db;
mem[481] = 144'hf327f9c303eff9bbf27000660d02ffcd086a;
mem[482] = 144'h0351f68f09720e940c57f7c1f26afbd7f1bf;
mem[483] = 144'hf4aaf8af0a5f0ebdf155fac200e7f8440e06;
mem[484] = 144'h066200e2f062f0300b8ffd7d04cd0256fd68;
mem[485] = 144'h081409c5f6b5011efe29038609100d3af5df;
mem[486] = 144'h0044081af146f6da03f9faccf5690bf9f730;
mem[487] = 144'hf2e20c7705820a65ff7b0640018cf347fcb7;
mem[488] = 144'h0109fbdc0ea9fd57f7f7fa72f76ef3a3ffae;
mem[489] = 144'hf61c0938ffa6f545f35c0384003cf5dcf8a2;
mem[490] = 144'hf68ff7d80855054b0ec2037403e70a5f04b3;
mem[491] = 144'hfa33ffa4f0a10334fe1003f20a6bff160962;
mem[492] = 144'h090f02e6f065f2bafee501b0effc090a009b;
mem[493] = 144'h097e09c006de081cfa8b0768070c03e60200;
mem[494] = 144'hf0d20eecf49f042efeec0e790133fa6efd79;
mem[495] = 144'h0b08fb03f984fcf2095dff7c0b45045307a3;
mem[496] = 144'hffa7fd31fd63fe480559f20e0e770e65018b;
mem[497] = 144'h031dfba3f97d0b690c84070af1a5fc68efff;
mem[498] = 144'h0a220ac30fe60053fc97f90301d2fcec0b59;
mem[499] = 144'hf257f95a09b206fe0e34077e0f36059f010b;
mem[500] = 144'h0a040a670719f07b0a77fa27f13e0988f4d3;
mem[501] = 144'hf4a5fcbd0f3c0bd9fe3afbb5f059fbb6fd57;
mem[502] = 144'h0bae0c080ca5f803f074f1b4f01afa5dff18;
mem[503] = 144'h066707790a5efa1508bc0b30f2b7f2e7021b;
mem[504] = 144'hf03607e00e23f025041e08b70eecf399fee2;
mem[505] = 144'h0189f094f1bf0ac704230fecfd68fbc2085d;
mem[506] = 144'hff4404d8fb3c008608acf032f6b0f749effb;
mem[507] = 144'hfb23ffe80ca3f15ef240f3da03b9fd1e0d21;
mem[508] = 144'hf07a0eed07bb069c037a041f0b32078df289;
mem[509] = 144'h0d7cfbbef88204a609aa04c9fdfbfb9dfb7b;
mem[510] = 144'h0b7a0d710fc801f30696078af2b803fef133;
mem[511] = 144'hf28bf247f1b80d67f04302cef638f0eeffda;
mem[512] = 144'h0ecb07ddf7da0de3f2f6f224f7620959f0ba;
mem[513] = 144'h072efe91f27a069e0b3a0ef2f77f0024eff2;
mem[514] = 144'h0a6e0b43f8d7020805830ceaf8a3fde8fc48;
mem[515] = 144'h01a3faeef0c304d8f5860f800c0400930578;
mem[516] = 144'h0bb402190be7f3110dfb0f1ff45204320126;
mem[517] = 144'hfb030252f8220f2c0f0f049ff3d701e5f66a;
mem[518] = 144'h04e00bb6f830f9a608bb061bf6b7f616f5fb;
mem[519] = 144'h08ec004a0eacfe170b05f29508ba03100408;
mem[520] = 144'h0efe079afc86f16e0306f1120edaf1000219;
mem[521] = 144'hff11f3c406d3febb0317f8d6f30ffc3107f4;
mem[522] = 144'h06f402d00a35f188f8f6ff42fdf70d56f859;
mem[523] = 144'h08a2ff9bf215fcd2fe360af90c09f3dd0689;
mem[524] = 144'hf46307edfd0f0f0ef09802b3fb3ff24c0a68;
mem[525] = 144'h013dfda0f44b0799f5470918f3af06a004ee;
mem[526] = 144'h0dca09380f4efc3c0f9afd35ffb2081bf8e4;
mem[527] = 144'h02fcf0c4f1340e4af0ee0be60f15022afbee;
mem[528] = 144'hfa8d09d50a6ff918f0adfe030043f70c0da6;
mem[529] = 144'h0382f4100b870a5002f0f1e2f39306e90b92;
mem[530] = 144'hffa400a906b80fcaf806067bf43705b2fcc3;
mem[531] = 144'h0f620bf6fbde0070fbb60656f528f271036d;
mem[532] = 144'h0c69f700fc65092ef125f843f7a00944f648;
mem[533] = 144'h0c97f8a9040902ee094d03af0492096ef43f;
mem[534] = 144'hf229f6bb01a5f407f029f0820117f8fc0d29;
mem[535] = 144'h05e5fed40421f5d7fcc60ee6f410048bf87b;
mem[536] = 144'h0c24fa9408e3007cf049f13409c4f1ca0455;
mem[537] = 144'hf266f930eff6010808bef95a08c2f634f966;
mem[538] = 144'hf138011c09950d0efb8efaf8f9f1fbbff76f;
mem[539] = 144'h05f305baf2c40a1c03d401a1f1f6fccf0f9b;
mem[540] = 144'h01e0062c0485fc9e0cb0f95f00d2fd40f8bc;
mem[541] = 144'h0ad306cef606053d02a1f63c065a06dffa12;
mem[542] = 144'h0276fc730b5cf8b2085d0d67fc250370f990;
mem[543] = 144'hf1b5f06df52104d80290fa810d8c09820bcd;
mem[544] = 144'h0cbbfd7c079ef6dd08820fe4ffcd0b1bf235;
mem[545] = 144'h063d0b0f0772f38d07980b3009190d6af277;
mem[546] = 144'h0857ff46054208aa0e650b4c0663fee1fa67;
mem[547] = 144'hf536f2fcffb10c0ff671f2c5fb4ef1c807fc;
mem[548] = 144'hf75ffa58f7e201b7f47802250b7ff1e707f7;
mem[549] = 144'hf469032e0063029ef68cfa950cd40cac09fd;
mem[550] = 144'h0d84fe0b036df51b0823fd50faef0e3bf9f4;
mem[551] = 144'h0629f0b2f0b2f83a01b4063af377f2160780;
mem[552] = 144'h0486085a0aa4ff3800f80fb00d7d08abf866;
mem[553] = 144'hf0ab0ca606c20f63fec50b88f82c0a7dff59;
mem[554] = 144'h041cf2c5f3590c860787f3ee0cc2f1340a62;
mem[555] = 144'hf6e3f724001cfa57f5bc081604ee03acf537;
mem[556] = 144'hf65ff7a9fcf0fe0af375f7a30a48092fff96;
mem[557] = 144'hf92df4cff8f2fd22f0fdfc930f2af1cef449;
mem[558] = 144'hfac8f557fe27ff70fc1a03a5063009bbf205;
mem[559] = 144'hfe5bf19b0e2b06c0fbc70375f504fd91080f;
mem[560] = 144'hf10a07e5f87eff150e7cfe4600cb0b3408a2;
mem[561] = 144'h007f0dcef0b903eefbd2f38d07e5f1ec079c;
mem[562] = 144'h0d480c79fd46fa0a03fdfc1eff8c0e8101c5;
mem[563] = 144'hf502f69dfee9f1ecf30fff10f1dbf8470f66;
mem[564] = 144'h040cf214f39307060736fb440d43fc7606e6;
mem[565] = 144'h0b3c0d38ffd50c410e5af54cfc540d93fa82;
mem[566] = 144'hf142f0b80a3ef8adfa990c34f54d0487f37a;
mem[567] = 144'hfa95fd99ffddf258008df26a02150e9dfbf5;
mem[568] = 144'hf2daf8980866f068009ef70b05d40735ffda;
mem[569] = 144'hf1a70039febef391f4acfa9ff1c9fb4afcc6;
mem[570] = 144'h093d0fa6f20cf3bcf733ff5b0bb804c30064;
mem[571] = 144'h0f3102e3f527fee20eb6070b0ee4033607a1;
mem[572] = 144'h0594fda90fec0a0ffe58fef20e380125f33f;
mem[573] = 144'h0ec2013ff3bcf3c0fcabf757fa520c960c3f;
mem[574] = 144'hf7baf9ffff360285f61901bf078f0f9fff27;
mem[575] = 144'h0b10f7f8fffc091f0ab1092e06480a72f9ef;
mem[576] = 144'h057b049500c3057efe10f60d0b790aaa0f63;
mem[577] = 144'h049202250853f771f17c04cffb55fbf70658;
mem[578] = 144'h0cd4f215fff1f1daf69f0441f5d8fb59f974;
mem[579] = 144'hf53cf9b0f155ff01fda40450fe36fe130749;
mem[580] = 144'hf7cefbee0b12f74f0be8f9fcf03efd670687;
mem[581] = 144'hff44024af7d30916f1a50e1f088dfd38ff2b;
mem[582] = 144'h0fb308b4015bfad3f31eefef0391f8d6fdd8;
mem[583] = 144'h0554f829f5b407cef91f0df10ec8f36b0888;
mem[584] = 144'h0485f5fdfc43fe860d47052f049a0c8e0b59;
mem[585] = 144'hfc650cfb06600427f6b9f685fb6bfda4fbe5;
mem[586] = 144'h0ef7f280f690fd960d00fdf8f26d0a2bfc0f;
mem[587] = 144'hf64e00d8f66d0e75fd8bf49cf29a0d01f56a;
mem[588] = 144'hf803027ffd4d0e55f4f1fcc6f49e0c87fbcb;
mem[589] = 144'hfa0c01e3f1bdf9d8fb1a0f2509580da3f33e;
mem[590] = 144'hf507f433fdb8fca5fd13f20dfb48f3d3f954;
mem[591] = 144'hf613006e0a68f841ffc90bfff93cfacf0518;
mem[592] = 144'hfea10db7061c0ee9fb1ef39205e0029a07d7;
mem[593] = 144'h0452f8d90437f218f944fcb60d2f06eff698;
mem[594] = 144'hf6db00210e39f164f382f0e1f33dfad7fbb7;
mem[595] = 144'hf282fb3e03c0f9f4f8bb00c8fe1df9180b70;
mem[596] = 144'hfe29f83d051af067fbf8f04cf7dd0535078f;
mem[597] = 144'h0d850f83f20e005ef09d00550c6bf664f1ef;
mem[598] = 144'h0660fce5f0d4f6aa0d170011f91ef9f30135;
mem[599] = 144'h0a40fba103aafc830d630eaffd8df01a07b3;
mem[600] = 144'hf259f12cfb18f0f2f571fe94ffe7f622060f;
mem[601] = 144'h0f12f8a5093ff4270bc1fecdf688fac2001d;
mem[602] = 144'hf068f2a5f8580361f0550578fd32fd7404a6;
mem[603] = 144'hfdfd0192030cf49c0c7604f3f533099cf885;
mem[604] = 144'hfd32fe2af2e80ac00acf0d5b0eb2f033f749;
mem[605] = 144'hf4e700a00712f43cf2d70f4cf2d30b68092a;
mem[606] = 144'h04d701180d43fc3b046f0a6f0f41f6fdff14;
mem[607] = 144'hf19d0b3afe9700750f36fa010f93f23a026e;
mem[608] = 144'h03990a98f90d05b8f31bf8aafd9300fbf9fc;
mem[609] = 144'hf08efae804050d4ffb59f4db0ea9fd590716;
mem[610] = 144'h015d03a70e7e09e501e40d6ff64d0c6efaf0;
mem[611] = 144'h06e307050243f5fff32af450fa69057c0f81;
mem[612] = 144'h08fcf85608f1f3d5f6eb05610378044d0502;
mem[613] = 144'h0152f059f5260197f6a80e47f232f652f29e;
mem[614] = 144'h0b5903b00ab9f24308af07e9f970fddaf16c;
mem[615] = 144'h0c32f548fbdf03b5fce4fc6fffbb042c0e32;
mem[616] = 144'hf95bfc8f0f1c085f031cf8970f81f9c70083;
mem[617] = 144'hfb710a7cf00b0ce00e2402b005a6f4aa0880;
mem[618] = 144'h0cc1f043ff69fbef08c005280ced0986f509;
mem[619] = 144'hfea20064f008f03c06fa01580499fa90f835;
mem[620] = 144'h033afb28018af903032ef0f30a27fc4eff55;
mem[621] = 144'hf5e40f0a0fd60667f2cc0faa0497f5b60301;
mem[622] = 144'hf6b4fb0cf143f31cf25ef1e3f62c03acf561;
mem[623] = 144'h087c030c08ce0808fc9af254f602fe8f0be4;
mem[624] = 144'h046c00f30bdf0c5e03a3f02ffd6cf2010784;
mem[625] = 144'h0728035007040afd0bf2088208effbe3fd19;
mem[626] = 144'h091c07790774fd2ef8aaff08f44f013e0407;
mem[627] = 144'hfe470c5cf964f4d5fff9f8cb0d420e2f0814;
mem[628] = 144'h06e8ff1efb790441026e0c570f7e0c540c83;
mem[629] = 144'h00bffe8b050d046cf96cfee7fb40f016fa29;
mem[630] = 144'hf5610f0f0ea40c29f423057dfff60c6801a0;
mem[631] = 144'h08f10740040bf4760cfb027109250b39f320;
mem[632] = 144'h03e2078e0989fdabf038f95a0729f768085f;
mem[633] = 144'h00c403acf7ce0d65f370f034f3e0f74bfc66;
mem[634] = 144'h0d940e85088ef7f40418f440f2e7f668024b;
mem[635] = 144'hf20103a805e6042d0fd2f14ef7b402cbf121;
mem[636] = 144'hf7580ac2fb460a36fadd07b10340f399ff6e;
mem[637] = 144'hf3f0f6f0f8a105ec006004610d20fa100d8b;
mem[638] = 144'hfbee0ef1f386019ff14cfdacf725f8ca0902;
mem[639] = 144'hf9acff0ff6b40aec013cf84efc2ff23a0854;
mem[640] = 144'h0502f76009da0214fbfaf7ff0d770b2ffb0b;
mem[641] = 144'hfaf2fca702f70a87f6740b32f970f51cfd37;
mem[642] = 144'hf630f75bfc4dfc2df21900a2fa4307be0509;
mem[643] = 144'h004cf1a7fdc10ca0f79c0f65ffce0888f470;
mem[644] = 144'hf7cef2fdf5e2f079f0d2fd7b0f53038bffb4;
mem[645] = 144'h0aefffe6065afa5afbaf0d9a0ec20f66fa0c;
mem[646] = 144'h060afc020a3bf4870e85f58500bafa2e02ad;
mem[647] = 144'hfeb2f9d80adffbabff4e0a210279fe15fa0c;
mem[648] = 144'hf0c40719f1f40e7709d40da1fc0ff04ff305;
mem[649] = 144'h07ec0284f2bc018a0008f2f3ffb103be0484;
mem[650] = 144'hf7ec01860fa3088cff34f7370d9ff9b9020b;
mem[651] = 144'h0eb505fafdf70b1c0c44f86708050551fc3a;
mem[652] = 144'h013a0ab3f9610f93f933050afa740714fef4;
mem[653] = 144'h0ca3f6480d00f100f9960913f231fd720a50;
mem[654] = 144'h067e0986f62ff9d7f07f0a970952fcf70fbf;
mem[655] = 144'h074b0271f45ff0e90666f3ec09dafceef96d;
mem[656] = 144'hf37af82805b8feeef1cff2f4f1790f2f0af3;
mem[657] = 144'h0754fc460efff1fcfa73f88f0402042c0ae4;
mem[658] = 144'h07e6f087f12a00bdf51208820e6af3f30faf;
mem[659] = 144'h035df24ff425f236fb0f093706ba042ffa3a;
mem[660] = 144'h077ff205f04b0e07f1640b7903c503b0fae5;
mem[661] = 144'hf58a069f0b3dfa840aff091d01b70d43faa1;
mem[662] = 144'h0aed060bfcaf0965faa10fa1f047fbbbf8a4;
mem[663] = 144'h090304c807eaf4a3fcf2f23efed10bc6efdf;
mem[664] = 144'hf4d8ff540520021802950b7af251f348fec3;
mem[665] = 144'hfb5903ac08e4fa6df98b06e404b508c4f9a3;
mem[666] = 144'h0ee0033bfb270ebdefd0f4150c1f0bd3fdd4;
mem[667] = 144'h0a560bf6f3720327f8680129f8d3f246f04a;
mem[668] = 144'hf52c0d9207ec074afffa05f307f00be40e4c;
mem[669] = 144'hf537f5e7f1910bd7040bf0effcbefca7eff8;
mem[670] = 144'h021004290c96f3c30b09fab1fb6b02c203dc;
mem[671] = 144'hf3230fb4fbb6098b029a0f64fa770d66fe52;
mem[672] = 144'h0e02f0d3f36bf7dafff508f80bd5f1e10802;
mem[673] = 144'hfc14fe6b0b31f68b018ff21bf863fa26f78e;
mem[674] = 144'hff37f47202a70c8cf195fac20107fe800e38;
mem[675] = 144'h0c42f076f9970eab01dd0ddd0544081df0eb;
mem[676] = 144'h0d0c0a20f2bf0ffc0dde0e550e580c110ece;
mem[677] = 144'hf8d60619f8a1f4bf0e22ffd10b2f08d504ed;
mem[678] = 144'hf758fe7900170e4803770c85f3c708d0fd63;
mem[679] = 144'hf8c50535fc03fb63065e0bb0ff230a36ffef;
mem[680] = 144'h0750f42e096b0bf0f90ff321077104b707c5;
mem[681] = 144'hf6e6fb80f0830d3708d4f19c0100f772fd33;
mem[682] = 144'h0099f068fc390130f25a012cf99802c6f88b;
mem[683] = 144'hf88efcf90dbbf74bf9a5f84afd1b02b9fb23;
mem[684] = 144'hfeafffeefb47f690ff6af1690b990ed408ce;
mem[685] = 144'hfbc0fb9c08b304d0f59ffa2f0b0ef334051d;
mem[686] = 144'h038ef060f3290f0df5cef617f552f5daf3d3;
mem[687] = 144'hf57bf34903e2f0f7005c0523fbfcfc57f849;
mem[688] = 144'h0fe209e9fde7f8b209160e9cfa70f579fd6c;
mem[689] = 144'hfd5005d00b8afb00fa0b0ad4f555fa83f637;
mem[690] = 144'h02a6086b01fefcfb05c00405f7e9f259fb33;
mem[691] = 144'hf3e0f5fc082806290152fae90a9c07c205fe;
mem[692] = 144'h0adaf21afa89fc1afcdafc09fbeb0886f3f8;
mem[693] = 144'hf4d60f88f07a0705f1d8f0330b05092ffd35;
mem[694] = 144'hf3c3fde9047afaab020f060af43804beff9d;
mem[695] = 144'hf1eb009a05c7ff310aa7f595faa0f5710ebf;
mem[696] = 144'h00cc05ba07890209f742f40e0033fb450c7c;
mem[697] = 144'hf03bfef50a76fda30718fa310e52f085f3a3;
mem[698] = 144'hf7a2015b0ef708cafe89f18bf02607f205fe;
mem[699] = 144'h0cef0328021a0ea70885fe92ff0aff58ffe8;
mem[700] = 144'hf8280629f32706ae0b67f786fe67f97bf4d1;
mem[701] = 144'h07b3ff3b08380edefbcbf2d0fedff88bf63e;
mem[702] = 144'hfba0fcb9f5190a2dfad50b0fff220bb9fa36;
mem[703] = 144'hf060f77b079201000df70766ff2cf12a0fc2;
mem[704] = 144'h04a7058f048c0172fab40615f34406bdf162;
mem[705] = 144'hf902f6ae0fa8f95807fa038700a1f3de0675;
mem[706] = 144'hf8560f07fb5c034908f2fa74fdfd0523f60f;
mem[707] = 144'hf949f0d4f0fff045fd4df68ff84002ad0e88;
mem[708] = 144'h0f0ff977f9a00ca5091ef681f74507fbf6ac;
mem[709] = 144'h0916f87d01a6fb96fce2f77a072501770a6c;
mem[710] = 144'hf197f79805eff18a0f37f30c0850effd034d;
mem[711] = 144'h0f4a020bf17401e4f5e50a8503e1f36ff08f;
mem[712] = 144'hf630f842ffc7fef7f2e3056000a00b41f2fd;
mem[713] = 144'h0549f9d6f1fe08daf858f942068f02a706c2;
mem[714] = 144'hf721001bfeb3f43102e0f82e0fdf080e0f02;
mem[715] = 144'h052cf78ff88703f605cdff88f063f6f300d4;
mem[716] = 144'hf896f75efa58f54ff9d00c1aff1cf0720101;
mem[717] = 144'hf9af02e303b7f6910a2603330d96fbd10be2;
mem[718] = 144'hf2ac07c2faa909880dc3f1d6fef60f310a63;
mem[719] = 144'h0fa409cdf151fa020480f6f2f01e0509f337;
mem[720] = 144'hfdd4f931f832f0d1f86cf387085e01e7f696;
mem[721] = 144'hfbe6fac40c4002f60e5c00c8f981f82b09d8;
mem[722] = 144'hf2b6fc4a0c25f30809d5f9e9056906840d6d;
mem[723] = 144'hf1feff00f89ff026fc3705c6089d08bc0754;
mem[724] = 144'hf4920922003502e1f7c3f5bb022af3aff4f5;
mem[725] = 144'h039a01a2f66103610e3cfe090e4506c30be4;
mem[726] = 144'h0476f57909310d9c0fd20c01f69ff2de0add;
mem[727] = 144'hfee608ca09c1023d0bb00ad4f403fe820001;
mem[728] = 144'h0d62fbba086303150104fd4d0a0fff6ef9c3;
mem[729] = 144'hf5ddf222f619f761089c0d7f0b29f4f800ba;
mem[730] = 144'hfe800984ffe1f9f6fd4cfe0c02a1f0e50cf9;
mem[731] = 144'hf54c0034f03ef64cf46b04e006230d33fcf0;
mem[732] = 144'h033cf14008c7f91c0f45f7b2f0fcf0820722;
mem[733] = 144'hfec90d0804d3f76100e5fd3206210fdff9d1;
mem[734] = 144'h0df4ff92fec8f194f874fb64f5050f000ed3;
mem[735] = 144'h0cee07440dd0f960f6d900d903c4ff59fc9d;
mem[736] = 144'hf108001a0a5bf6b4f0710c8df6ae07740af5;
mem[737] = 144'h0550064e05920f030e7bf7d000190d6c0673;
mem[738] = 144'hf98a0fca03f7fac0f87904ac01860d68f93c;
mem[739] = 144'hf497f7c80fde0b4afc01fb51fd23fc8d077f;
mem[740] = 144'h0b6bfe9afc5f0ab80379f9cd01ecf68709d7;
mem[741] = 144'h0426f1b10d38f007f6ea0c35064af1f1017b;
mem[742] = 144'hf26e04730be508a3fe790cec0016f7c20c78;
mem[743] = 144'hf4970dcc06fc09690394002901aa0da8fd21;
mem[744] = 144'hf6c30ebd01db0dc4f43c00380a9ef4e6f3dd;
mem[745] = 144'h00f5f78cf23cf7b40ab6063afeaff41efc2e;
mem[746] = 144'h0f0c0049f537f6c90678f678f8cf046a0552;
mem[747] = 144'h08ef0b2efad30593f916fb920226f0c5f487;
mem[748] = 144'h07cbf7b0f322f62f010a0a820b76f3c1f296;
mem[749] = 144'hf1a5f28d0749039af7da05b7f644fd8df30d;
mem[750] = 144'h0a9707b80605fef00986011efa00f00cf44e;
mem[751] = 144'hfb62f186070702770a64f8c60b2308aa0672;
mem[752] = 144'h0fde0b25008b0d0df34c0eca0811f1460c5c;
mem[753] = 144'h0df70d5603cff76e0f65f86ff338f8b8fc1f;
mem[754] = 144'h0d59fa7103f7f4a20cabfde0037d051f01a0;
mem[755] = 144'hf22c0d6ffe4dfef3f8fbfe07f1c7035ef596;
mem[756] = 144'h08620d200dfeff6f0c940b35f8fef3b8f227;
mem[757] = 144'h0766f80cf8cdf471f1830d39f226f1f9fad1;
mem[758] = 144'h08a9f067f75bf7f5fc090cfef77af85fff92;
mem[759] = 144'hfbed0ed2f1230a26fe2600a30d5f04c10a78;
mem[760] = 144'hfb4af01b08c0f067088df0270e4cfa58fffc;
mem[761] = 144'hf86a03630806f1f5fce2f3370a9f0345001b;
mem[762] = 144'hf4250840f1e20766063a0c5f0237062c02c6;
mem[763] = 144'hf5a4f1d509fef4dbf03efdf50dc6fce10b49;
mem[764] = 144'hfbfdfc9efa77f2b7ffcafcb7feedf786f3da;
mem[765] = 144'hf5330a02f6f7fcb8f706fb330154f89ef2d5;
mem[766] = 144'h0d8808b3fc6905150549f6b0f1850c5dfa1c;
mem[767] = 144'h044508690f03f7c5fb9f0a48fcebfb20f779;
mem[768] = 144'hf5d0ff680ffa0ceb04d8fcaff32f0d230cf3;
mem[769] = 144'hf17605f70d4afe62069f0ba901a00725f54a;
mem[770] = 144'hff0ef463f976f7d60374f34a0b9e06150d6b;
mem[771] = 144'hf5ec06e8f4e30ac6f5c10d140bdcf7eafb5f;
mem[772] = 144'h0854019ff51af1e6042400d10be90aedffb3;
mem[773] = 144'hf3c90138f7530edbf03b03f4f94803670157;
mem[774] = 144'h01d4f059098b0103f10102240530f399f7f7;
mem[775] = 144'hfce9f071000e003104edfbbdfacbf0f906ff;
mem[776] = 144'hf510fd7c0404f8fef17b090dff9102f6085f;
mem[777] = 144'hfa76fdd3f4ab011b0e17f83901aa0712f245;
mem[778] = 144'hf5280f53ffbf0b2f03c20254011cf76efd72;
mem[779] = 144'hfca70608fbe8f2faf73cfd81f9d30cf60bb3;
mem[780] = 144'h0ddcf8bd08b9f7ea0738fc1c0007f169013d;
mem[781] = 144'h0563febff5ca01340beff013f635f15bfb83;
mem[782] = 144'hfb0705d70bc4053406160fd0f8680990f3af;
mem[783] = 144'hfb5ff928009c0a2c0909f2dffe5008c40525;
mem[784] = 144'hf645fb88f566ff1c0f870b50f237fee5fbdd;
mem[785] = 144'hf3b0045f0d08f7a2035df81bf0320abef7fd;
mem[786] = 144'hf89ffc4ff263fc20f075f78efc2e0b51f2e1;
mem[787] = 144'h0899ffa20c5bf70ef4120aac0f1df9490263;
mem[788] = 144'hfeb3fdbc08f3febb0d920a820b0ffc350326;
mem[789] = 144'h0f2aff9a0091070ef708ff03f64ff7e5f805;
mem[790] = 144'hf302fd350810f2570701fd100489ffd4f4d8;
mem[791] = 144'h01dff12d0daf0019f3ca0d8efa7c0fd4f156;
mem[792] = 144'hfbd7087509adf26bf065f065f5c40cc20552;
mem[793] = 144'h0f4bfde8fc79ff96f07ff6e8fba207820312;
mem[794] = 144'hf0470d39f546fff7fd160373f87df94b0134;
mem[795] = 144'hfd4bf7ec0ae8fc95f7cb0885f103f4d5f1a4;
mem[796] = 144'h080df3b7f9d4f66df5e2f53b08a50e82068f;
mem[797] = 144'hfac5f303fde9fc51f45e0fedf878f068f3c9;
mem[798] = 144'hfb11f480fb350a750f26f928050407c3009a;
mem[799] = 144'hf47e001df2f70bc2f67df881f4b50292f123;
mem[800] = 144'h0f28014cf4d8f3fafbce01fcfee9f2fcfaa4;
mem[801] = 144'hf9ef0701069d0fd202ac0dfef9c7f4ce0ce6;
mem[802] = 144'h086a0201f966f8a3faf60f1807f7fef8f839;
mem[803] = 144'h0cb9f27ef0de0997f055fc5df3bef09efeab;
mem[804] = 144'hfc4afcbef5a7fa320fddf36b04bcfe80fbad;
mem[805] = 144'hf3f7f99df7fb0d0f05510a24f509efd5fb8e;
mem[806] = 144'h0749fa1f0f330afbf7d4f2fd0b30feeb03b0;
mem[807] = 144'h09350e51f7b40664068d062f023a020e083c;
mem[808] = 144'h0779fa670139052f0a290594f5a907cd03a7;
mem[809] = 144'hf626f2cffe75095e036bfa35056f0c11041b;
mem[810] = 144'h0537fa63093e054afb6a00ca0093f691fc03;
mem[811] = 144'hf6a2f3c80ceaf1f10e450e7b014efa6e0e61;
mem[812] = 144'hfac9ff79f5ecf8e90c56001e0b840756fbb3;
mem[813] = 144'h0aeef418f2b5f815f0520df60ecdf0470077;
mem[814] = 144'hf9630725073202f603580bc4fd1801a2fc6d;
mem[815] = 144'h0933f631fc640ea3f0fdf4c105d504350d03;
mem[816] = 144'h03e5fcedf085f25c0f0af3be0d3c0f6a0561;
mem[817] = 144'hf5e4fb99fe490963021c0bbb0ea9f039fe17;
mem[818] = 144'h08b50448f782f6e60113065df503feabfdaa;
mem[819] = 144'h009500f6f3b6f7f40819077c0044fb1d0aad;
mem[820] = 144'hf370f20609c40d20f4cd03bf0728f25d0608;
mem[821] = 144'h0cdaf482f084074af438fb9af97908840b30;
mem[822] = 144'hfd71fb07f38e080afd0401670bf601270b7a;
mem[823] = 144'hf885fbf30d79012af34b0fb406050a16f5db;
mem[824] = 144'hf0f5f04ef7f904180ab50cbf0320070bf610;
mem[825] = 144'h09aef1e6f65e05abf514fb4508800b20fae6;
mem[826] = 144'hf4b10195f80afdc3f06a04930bb60afbf3ca;
mem[827] = 144'h0165f33902ee0897f171069d00aafe08fbbd;
mem[828] = 144'h091209bb0da10e8b05c6f4a6f34efeb8f316;
mem[829] = 144'h071bf6d1088105bf064802a5f825f332031e;
mem[830] = 144'h063701b2f04f01a5f64ffbd3f89700c30505;
mem[831] = 144'hf4c20a34f0a10730fb430fa40e8f0ad609da;
mem[832] = 144'hf38df25e0238ff26f46a0137003e01c4f296;
mem[833] = 144'hf2f10422ff7a0b0aff55f707fe7b0a5afbc3;
mem[834] = 144'hf0ae0154fb1104470416051af1dc09cb027c;
mem[835] = 144'h0b070550f8040ff10021f94d082df4880a16;
mem[836] = 144'hfe9306eb01ff0cbbf0cb0223f889f0ce0b6b;
mem[837] = 144'hf288faee0f25ffed06810545f83afd8e0b96;
mem[838] = 144'h055cf7ad06c9f59d0a51fdec0e420db70c6d;
mem[839] = 144'hfb9e02b0f4d10cf802260f010408fa190310;
mem[840] = 144'h01f10c3c0c90f2edf5910ec30f05f437fd82;
mem[841] = 144'hfea30becfa450652fc280b03fec4f8b9f735;
mem[842] = 144'hf66a0b21f5eaf7370ee1f9510f16f3080f05;
mem[843] = 144'hfb76023b038ff7250a2f08580912f0b90fec;
mem[844] = 144'hf69d0efb0233fbc7f3d8fb3300f1016d043f;
mem[845] = 144'h0f07f7ccfe1b0703011efbfef1ce043b02ac;
mem[846] = 144'h0842007cfec9fc140d36fc6b0039fb3604e1;
mem[847] = 144'hf8ea0fc1faf006cc0eca03e00a10020a0cd8;
mem[848] = 144'h013a070b0983f08d08470acf0eafffa9fd71;
mem[849] = 144'hf1b7055bfaed090df839f180fdcc01660901;
mem[850] = 144'h0c28fa130b260997fe4bfa6ffade0a640cc8;
mem[851] = 144'hf751036a084b0df90700f943f385fd2bfa5c;
mem[852] = 144'hf4b60709ff0a04d60d29f859f3e70ec10cd2;
mem[853] = 144'h0bed0aa70c8d0434fc1bfaf4f6e00f83f22e;
mem[854] = 144'h09b2fce6051a0a3601e803fd09ccf1c9f4d3;
mem[855] = 144'hf3ad023af7260e2c076df2d40d94f36602f9;
mem[856] = 144'hf6cf0c800b220530090af75c0d8d08a20e5a;
mem[857] = 144'h0221f51b0e72fb2ffd63f34b038dff91fb81;
mem[858] = 144'hf8bb0717f9cbf989f475fa630bcaf61a0834;
mem[859] = 144'hf1f9069303380cef099e0908052af6730146;
mem[860] = 144'h08c9fc8cf69bf7230530f0140fd6071c0053;
mem[861] = 144'h01a3f7a4f3e3f8acf652fc81fa5af159f78a;
mem[862] = 144'hf36408ae0d98f2290388f6e7f881fb9c034d;
mem[863] = 144'hf9030a1b0510fd51f727fe430eb00ad1f0a1;
mem[864] = 144'hfc97fc83f18b050208340192faaff46f0ad9;
mem[865] = 144'hfe20f31f02faf961fd810d09058f0d9a016f;
mem[866] = 144'h098af519f521f6ac09f4f0a20a26f618f6fb;
mem[867] = 144'hfdb5fd6c0cbe01b9085af97ff115f4e5fec6;
mem[868] = 144'hf96507b7fb81f7dff4bcf012f4d3f5110e72;
mem[869] = 144'h035b04280eb1ff82fb96f3f500d5f23f0e3d;
mem[870] = 144'h0c79f18af5dff1140279f6ddf274f2b20335;
mem[871] = 144'h008cfd320abf03280d68fbdbfa9af1e00b1d;
mem[872] = 144'h0d61f29402d7f377f9d5fc3f01b9030df452;
mem[873] = 144'hf5f2f487f50e01c705ccf474f63ffbdaf12f;
mem[874] = 144'hf6ef07740c020fd5f7090993f1af086b01fe;
mem[875] = 144'hf14902000d11f70bf9c7f3c00f8f0f5a09c4;
mem[876] = 144'h0830f425f66a092a09def82906acf0e8f5c7;
mem[877] = 144'hfd0eff61f909f0a1f0d801fc06e50d1e047a;
mem[878] = 144'h0933f7cd0800f1fbf51cf8700912fccbfa08;
mem[879] = 144'h07f702a90e800acdf58df3ca0073018a0ca9;
mem[880] = 144'h06a40402f8b40810fe80fe39fde8ff57f2a2;
mem[881] = 144'hfdc4f703f7550efb00710b70f815f292fd33;
mem[882] = 144'hfa5ff4c7f50c0caef4a2023dfc13f0d10ef1;
mem[883] = 144'hfbc9f377f70f0d2af87bf09afe1d0a850570;
mem[884] = 144'hfc28060ffbe5f77df2e0f931055e0de00ccd;
mem[885] = 144'h0b15f7c90ad2fcf70e99feb7fa24f3caf047;
mem[886] = 144'h053a0e23fb1ff059f9800440f97709720a7b;
mem[887] = 144'h094e00cf08e407110bef00cffd260bea0b4b;
mem[888] = 144'h006207b7f179040b0d95024bf9110f7801b4;
mem[889] = 144'hf3ab04cd06b000c5fc27f66105710849f58b;
mem[890] = 144'h02cd0dfcf2e70a33f9ea08e7f774f6cc0d4e;
mem[891] = 144'hf7fff2aa0a8600defb1c0b3005f1f36408f7;
mem[892] = 144'hfa2a0884fa1cfce20265febf06bdf0620889;
mem[893] = 144'hfc32f0f80223059f0ca90f29f168fc6cf02e;
mem[894] = 144'hf87a030d08f307a5fb320b42f4a20a57fc6e;
mem[895] = 144'hf39b0c70f517f0320550fe75f92401380b93;
mem[896] = 144'hfa9aff66fb3cf444f9510d8ff7fd0c49f6b8;
mem[897] = 144'hf026f5230e510f8d07f201ebfa68fb59fe6c;
mem[898] = 144'h0566f454003e07dc0f2df1270f1df1cbfde2;
mem[899] = 144'h063f0a0705750439f5ff0d4ff426079e02ff;
mem[900] = 144'h0d90f850fc3f018c06e60a47fabff791f035;
mem[901] = 144'h06e2ff48fc1cf88af292f130f9190edbf24f;
mem[902] = 144'h0a64f0f8fc3f069ef9030ee4f340001409a9;
mem[903] = 144'h0cb9fbd4065efd9cfba5f25cfa93f249f4bb;
mem[904] = 144'hf4f3f075ffbdf55d0bfb0a04f709f046f14b;
mem[905] = 144'hf83df2b5f766fc11f7e7f155f61b0988f38e;
mem[906] = 144'hf47d0562042ef9ef0c5804110f73f170f4e0;
mem[907] = 144'h0716f7a50a73fad9fd9e061f016f012e0519;
mem[908] = 144'h0116f39b0c17f91d02010444059a0790fa3b;
mem[909] = 144'hf64207050e92fd8a0e000438011cf93f0c3d;
mem[910] = 144'h0060f4b0026508a10384f06afdc909a5f885;
mem[911] = 144'h0f3806d9fa6b00b5f05504e606d70d3bfbbc;
mem[912] = 144'hf4a7fb1b0581f45303850f9c0f5107d10b9b;
mem[913] = 144'h09a3f669f64cf67ef882fca8f079f68d07e8;
mem[914] = 144'hf97a06a7034801180a8cf874035cf48a0900;
mem[915] = 144'h0e37f7ea09f708b9f20105ba0f15f2f9f40d;
mem[916] = 144'hf605f014f82bfc77f5990ca4039af24ef155;
mem[917] = 144'h0eb50fc3f2a60c0cf823013ff2620c0007e2;
mem[918] = 144'h0ec700c502360cf5f8840601064ffc1708bb;
mem[919] = 144'hf4470ac00af6f02506740651f75ffff00776;
mem[920] = 144'h0a61f27c07f1f98ff6770be6084b0a5cf5f4;
mem[921] = 144'h03ab08c709bb07c70890021801e2028405eb;
mem[922] = 144'hf9d5ff7ff5000dbef370fe5dfe33f59ffab7;
mem[923] = 144'h0adc0435fe8fffc00a4f0f8303e40198f2df;
mem[924] = 144'hff0203af06cefd42f832fd980316fa72f2fb;
mem[925] = 144'hfde20b6e0572fac90f3b08f10281ff810168;
mem[926] = 144'hf8ea01d80f56f65ef2e506ba038403cbf2d3;
mem[927] = 144'hfed40502f0920afc07ea0d310d6cf1dffefd;
mem[928] = 144'h0b34ffd80c7308b0f9a7fe70023808f50a2c;
mem[929] = 144'hf7fc0b59f09005b4f296ff1c0d5a0464f08a;
mem[930] = 144'h0d9efea4f5200efffab7f617fac4f54b00b8;
mem[931] = 144'hf6de00120e570218fd64f77a0e120a18f07a;
mem[932] = 144'h04f3fb310f1a0827f51c0fdd08cb05800bde;
mem[933] = 144'hf630073107650ce6fd290ec30c27f7a4fbdc;
mem[934] = 144'h07c400adf647018806820c48fe42f3930c04;
mem[935] = 144'hf736027af3ed00c6fc2bfb16fcc0f5730b9a;
mem[936] = 144'h07fff8d70ca0faa0013df533f6c0f47b003c;
mem[937] = 144'hffe200a0090505b4f5c90b230e5d05b60720;
mem[938] = 144'hffa4fac0f293065ef515f056f918fdc3ff1d;
mem[939] = 144'h08c60e51f425f8d405100c260ed9020cf408;
mem[940] = 144'hff72032500d1049a0c260d3ffddbf4a80cc8;
mem[941] = 144'hf917f5c0003bf30ef3420e09f360fdf0fd15;
mem[942] = 144'hf45201ae0b79f12c0b51f59a08270fa2f249;
mem[943] = 144'hfb3cf54e0a2e0329f5d0f228ffd3f43e0705;
mem[944] = 144'h02a2fc04fb67f18103cdfd660ef40d420243;
mem[945] = 144'hf23401c00067fddc040c0356fc13030500f1;
mem[946] = 144'hf905f395043c020903b5fe5b0db203f1fa85;
mem[947] = 144'h0818098b0bbef614063bffb70ddcf71cf3c4;
mem[948] = 144'hfc820cad0522fc8cff53f045076ef2affe33;
mem[949] = 144'hf22bf0b2059bfe950646f5acf42b0046f677;
mem[950] = 144'h025cf270f5250a3ef74a0d61faf404affc8c;
mem[951] = 144'hf994f393f4eef6a3fe04f35b0e4af2ad0e25;
mem[952] = 144'hfac30569f26e0ae807190140fe010e01fd4e;
mem[953] = 144'h0f63f784078902b40fb4f9f00e8ff6f4efc6;
mem[954] = 144'hf03e0ba108280b5af177f3df02720648f877;
mem[955] = 144'h09ad0646059ef494f4ee0bbff3c50cbdfdbf;
mem[956] = 144'hf303f76df1d8f53807c10746f494f7750658;
mem[957] = 144'h08890ee90738f6f501c0f4200e1af19b062c;
mem[958] = 144'h03aff46ff0de040cf3aefb8efe4df5a50537;
mem[959] = 144'hf285fc59fa0903f707db073e03f2f7aaf47d;
mem[960] = 144'h09bc03370ea0fc3cf3e202f9fd5ef701f19e;
mem[961] = 144'h0d7dfdc4f97bf7c7fe2f0521fdaf0c6bfcb1;
mem[962] = 144'hf567066c0b01f6f4f9b508960cbff0eefdc7;
mem[963] = 144'h00a2004afc8c0cee0f3a093b0f7af369f71b;
mem[964] = 144'hf62d07c7002bf87e0e5c0773078df1fdfe29;
mem[965] = 144'hf2b101a9fdd5fd5007e3f13e054ff2770aab;
mem[966] = 144'h0e72f74c0d2bfb3a01c10e1809bef8420a9c;
mem[967] = 144'h001106e6f665f5caf75a0e24f622f28bfc25;
mem[968] = 144'h03d3fa1b0022f6f00982f0ebfb31fad80d90;
mem[969] = 144'hf484f40b07abf230fa38f07b08ecf6ad052a;
mem[970] = 144'h015ffae9010af37a09bc082e0ce3fdf30be6;
mem[971] = 144'h0e42fcd8f2a2f9310a940e90fa2bfb9408f4;
mem[972] = 144'hf969fa05f1ba0be2f7fb0d6ffb4f02e8fb7b;
mem[973] = 144'hfc91fa7902a4f338fdf104e106810c66fead;
mem[974] = 144'hfee8033cf918027a00780ab4ffb2023605af;
mem[975] = 144'hf03d012b00a4fb1f060306f201730d23fd0f;
mem[976] = 144'hfbdff4780fe5f7990fc1fad5f5e502defc3d;
mem[977] = 144'h08cdfe280c68fdb3001cfca5fca1fd79f7c7;
mem[978] = 144'h07d8f5c209070b72f2da04180b38ff1a06f9;
mem[979] = 144'h0852f9af0dfb00790192fc2a062d0535fe5f;
mem[980] = 144'hf103f965f656fb1907b6f2b5f1e9063efa94;
mem[981] = 144'h0ec00470f4920176f11dfe42f00a04510b52;
mem[982] = 144'hf6dffc45fb55f9b1fa650092f1ce00a703f1;
mem[983] = 144'hf70cf2cc01070e7a029af6990376f821f2e9;
mem[984] = 144'h0390f150f08809f80b2d030dfd780358035e;
mem[985] = 144'hfb51f3e3f2b8f49ff3d7fd7108af05ef0e4a;
mem[986] = 144'hfc85fb1906a8f7640a3ffe20fce9faa3fdb7;
mem[987] = 144'hf7b4f4ddf1d3f2260bf0fb1afb9b0d94f88f;
mem[988] = 144'hf4cf0cdcfe0e06d9f4d103fcf69a0992ff04;
mem[989] = 144'h0fd6f0bff04800b9013507fafe430fb4fe51;
mem[990] = 144'h01080733f1580e4cf64e0ad7fe0707340ce4;
mem[991] = 144'h001c0567ff12f7c1f780025706c2febe079b;
mem[992] = 144'h04a20331ffaa0eb4fbc3fe02f8840cc3f166;
mem[993] = 144'hfe9bf460072307ba08b7025ef002f946f517;
mem[994] = 144'hff2b0992f86e0b8f00abfa0df82605b10d4f;
mem[995] = 144'h0c170b84fdfa0fbcf129f6f906720e880118;
mem[996] = 144'h09a5f5cbf3350de505830444f741eff70df2;
mem[997] = 144'h0ed3fc10f9cb090c08befca40c610382087e;
mem[998] = 144'hf66dfd88f1f104ecf88af5b1f5def0fef657;
mem[999] = 144'hfbbbf8610bdc07a6f03bf014f4bc02aef621;
mem[1000] = 144'h0373054bf61601f6fed40c6f09aff1f8fbe3;
mem[1001] = 144'h00b1f155f999fa07089d05f0ffbd0c3f0501;
mem[1002] = 144'h0179f6f6f3b6ff2dfb1806b3fe8bff870803;
mem[1003] = 144'hf291f4b805d501bcf3d5fae906c7fd19fa46;
mem[1004] = 144'h001c00a1017ff51a013cf304f6700365f61f;
mem[1005] = 144'hff7d010efc75efc9082e08cf04e1f4560bd2;
mem[1006] = 144'hfe030e4503e309e8f36b0fbcff2df1d4f6da;
mem[1007] = 144'hfe65085d08a60b7502aef17705c6ffb8febc;
mem[1008] = 144'hffe00922008ffc93030cf2450e4cf9adfcbc;
mem[1009] = 144'h053df4b50fa2f2310ca1041a02ee00c6fe8f;
mem[1010] = 144'h04e90072fa12fa060a68f958f922f3a30c78;
mem[1011] = 144'hf799f1bdf50afc0902a006fbfbe109e60f81;
mem[1012] = 144'hfa02f5360c6dfbf6f24009c3feebf50406cf;
mem[1013] = 144'h0dd5f7f3058df1ddfa100ed2ffe105a4fb06;
mem[1014] = 144'h0f5d0886f611f19af8480a12f8cb0e92fbd0;
mem[1015] = 144'hfc06f303029af7acfcdc0ba8f7fef8bffb8c;
mem[1016] = 144'h02d90228fbc502ae0b74ff30f0c2093ff1bc;
mem[1017] = 144'h05c50911fe700be10ea4f47bf35cf7e9f09c;
mem[1018] = 144'h04d5f228fc1c0d3d0fc40ea9f049f0400c43;
mem[1019] = 144'hf6d604dc00a00157f3250c22095208170d43;
mem[1020] = 144'h036b09d9f0cff2990a7807c6064dfc740ba9;
mem[1021] = 144'hfee7fa57004df6a1fc9ef290fc29064b0f1f;
mem[1022] = 144'h09a209e304db040dfc2104c2fd640c84fb27;
mem[1023] = 144'h0e15f8e6fe77f6f4f82d07f1f43cf1240529;
mem[1024] = 144'h0fa70746064108ec0ecaf5bbf225fbdff8b2;
mem[1025] = 144'hf9b608b7052c0ccdf8c8fdb6f4d9ff4c079f;
mem[1026] = 144'h0eee0170f5dbfa76086ef27d08f4f756f448;
mem[1027] = 144'h0e110755f9e9f698f8c008b1f20d03d206dc;
mem[1028] = 144'h07e6f26cfb9dff70f9cb0a8f0cc4f8c90e0b;
mem[1029] = 144'h05d901a9fff8feebfd2f05690ded0ad50ef4;
mem[1030] = 144'h005e0b300022faac000ef17707fa0db606bb;
mem[1031] = 144'h078cfc95fa54f342fc4105b50995f7750d92;
mem[1032] = 144'hf0e1f59d0731054e0438f85ff754f8da016c;
mem[1033] = 144'h007ef258014c094afc83f7cd0d460b11f19c;
mem[1034] = 144'hf2410dc802950329f8b1f7fc0f6df182f747;
mem[1035] = 144'h0f3ff1160d66f09a0618001bf7cf0fa0ff70;
mem[1036] = 144'hfdc102ac058bf3d0f748f2eef59402870cba;
mem[1037] = 144'hf6f8f802f126fb09f9c7fa5af53305e10315;
mem[1038] = 144'h051dfda8015f0f8d0eb7f977f8c3fa65f578;
mem[1039] = 144'hf20f0fc4043a065cfe9b00c8070d0c3300ba;
mem[1040] = 144'h06fafb930556fe27f1e10f030f6502a4ffc7;
mem[1041] = 144'h03400f220542fba4f1fcf5dc0f19f7d40d94;
mem[1042] = 144'hf9f7f684fe4c0adf0e4ff57e0670f93df3d3;
mem[1043] = 144'hf0d60cc205c1071f0150060efe2ffa7e0f51;
mem[1044] = 144'h02e2fdc7fe73f79e0dfa02260165fa0200fa;
mem[1045] = 144'hf46a0823077c088df2ca073cf079087afa31;
mem[1046] = 144'hf77b0e2efc7d0bfb0215f419fcec0097f0b2;
mem[1047] = 144'h09ea04cd05ec0ff6f488f573f75df687fdfc;
mem[1048] = 144'hfc5900e3046cf538f709f5bc0cdbf0e400b1;
mem[1049] = 144'hf2e4fec2fd9305510599f6660b48f3d9fd4b;
mem[1050] = 144'h09daf98c03d6f81dff78f3840cc2fb6b09ae;
mem[1051] = 144'h0d27fc78fe660b7df1c70a16f7fffd93f67a;
mem[1052] = 144'h0a6ffaa007790fa9f2e3fde8ff06f15e0ef7;
mem[1053] = 144'h01f6f238ff76f10601790149017f0d97038c;
mem[1054] = 144'h0fdafc9ef090fe360130f133fb7801b40bf7;
mem[1055] = 144'hf1360f410a03feb503d9f1b50363fd23f3ab;
mem[1056] = 144'h04960c3e03130ebd022f01b40ebd0e040f17;
mem[1057] = 144'h0561fdb4f55800fe0d97090d04f40e640d1e;
mem[1058] = 144'hf25008e6fa71ffc1fa8f0711ffa3f5620c8b;
mem[1059] = 144'h01dafeab0de2f9fcfdf503c0015af8d6f1b4;
mem[1060] = 144'hf97cf8b1f21200ff0b6cf852f1d406d9f0b2;
mem[1061] = 144'h04baf30204af0689fb0af368061ef18501f5;
mem[1062] = 144'hfc23f3b40ce8fd13f3cd0dbcf9fb03f9f903;
mem[1063] = 144'h08080e32f25a050d07abf5a4fbcdfa17fc00;
mem[1064] = 144'h0e2d0e5d0f5afe6ff4510bc00ab50a170c92;
mem[1065] = 144'h0eaf0b3ef71efccdf95bf874f6170445f483;
mem[1066] = 144'hf2130d44f828fe0808d5fc45fe6b086c0e99;
mem[1067] = 144'h043605db091dfd1dfc1d0af70efc02ff0c08;
mem[1068] = 144'hf775f1bd0e2303a4f72f0f6a0a9900e50938;
mem[1069] = 144'hff47f2bd0dc00e76fd1902460c10f8ff05f7;
mem[1070] = 144'hfd9afad7f8430e4805c201df02510d72fa11;
mem[1071] = 144'hf8ea0c31fdaef737033c05990597f7720c5a;
mem[1072] = 144'h0a6a0469fc78fea70ecdfed3f05cf00f02e0;
mem[1073] = 144'h0ea1000305fe0c210b0700c50134f6a2f0b8;
mem[1074] = 144'h095300d9f8f4f1a9fc78f2dc0ef7fa5b04e6;
mem[1075] = 144'h0c7eff050e51f3c3f3c008640149fde60461;
mem[1076] = 144'h0a18f7960b39f6b90c81091a096c024c0a40;
mem[1077] = 144'hfd0afd4ff2200594f418ffd008e7f296f706;
mem[1078] = 144'hf6cef5edf7a5fff1f173f8f3fe080afe03d0;
mem[1079] = 144'hf66ff7f5f928fefefa5a0ca1fa1e0e05ff18;
mem[1080] = 144'h05130e59fc54fb73f49a0d520a9a08b70767;
mem[1081] = 144'hfe3704d5fb500e6ef7410430fc140e4afa90;
mem[1082] = 144'hf361f7150817f540f524f7faf01103a8f537;
mem[1083] = 144'h0fb90e70fc14f745f8df035e0f0bf42a03fd;
mem[1084] = 144'hf652f47c0468f88e0fae0c910b5cf026099b;
mem[1085] = 144'h05c10054f71405df00e50c18fc53fe64eff3;
mem[1086] = 144'hf9e90228f6b4ff2b0d8f05bb05e6fc05fdc8;
mem[1087] = 144'h00ac0c1107f10ad2f9d1f19800dfff050e54;
mem[1088] = 144'hfc0dfe02fc45f8cf06fafc5a0e740c32f265;
mem[1089] = 144'h0c2e0febf6ea01db02920eeffb1900f10c03;
mem[1090] = 144'hf464fafafd98fbd0fa78033a0746f2af03b1;
mem[1091] = 144'h0c0af7ab074a0abd0b3b03e7002b0dbcf2b9;
mem[1092] = 144'h01c60e31007202cdf7aeffd8fa08f83bf1cc;
mem[1093] = 144'h06b80f7c1078fb9c0008f02ef2770fa60922;
mem[1094] = 144'h01a6fbedf9de02d0090f084e01b300620c16;
mem[1095] = 144'hfa5f0b14064a0ccd0a68fd7d08a9fa1effed;
mem[1096] = 144'h0d370f2f0ac0fda3f573fd83fe9502d0f2d6;
mem[1097] = 144'hfc4e0a110e15f2cd08a6f7fc07d5074a0b87;
mem[1098] = 144'hf3baf36ffbee03a10d0bf23601b1f60103cd;
mem[1099] = 144'hff93f76f08b4f3fc07d6fd2b0d3afc3f018e;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule