`timescale 1ns/1ns

module wt_fc1_mem2 #(parameter ADDR_WIDTH = 10, DATA_WIDTH = 144, DEPTH = 1024) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'hf5d2f5ee00a3fc4e05e30c82fbae023c0dbd;
mem[1] = 144'h02adfcc6f81a094a04dff0fdf555f4d70308;
mem[2] = 144'h0169fdaaf83bf5e30dd00d230c8df4a8f8ed;
mem[3] = 144'h0d5b004d0539f1fd06a1fdc4066effc80f93;
mem[4] = 144'h01f2fec9fd55fe3cf1f109d8f978f32cf70e;
mem[5] = 144'h09b20d9a0f520368f028040ef155f99d02a9;
mem[6] = 144'h0075f894099df25af198f4450da2f2cdf3bd;
mem[7] = 144'hf97afd350198073f094f0231fa20095bf27c;
mem[8] = 144'hf4ad07b5f601014a01df0b7b0f61fe400ef0;
mem[9] = 144'h011200c1f53b0e1d0361f790027bfd44fceb;
mem[10] = 144'hfc13f58e0ce7048dfe44f507f3c706cafd07;
mem[11] = 144'h0f0b025403cff0d50406fe68fffa02b10786;
mem[12] = 144'h0970f3a3041ef13af66d0adbf575f38bf969;
mem[13] = 144'h031e034df1cfff360e72f769f443053a018f;
mem[14] = 144'hff660047fca70f6af9b0fde6f19ff6ff066d;
mem[15] = 144'h0db0f7fff4470019f141062ef0aafc820232;
mem[16] = 144'hf218f953f7370bf301bf02c102b9fd81fcca;
mem[17] = 144'hf9fefbeff53500c702440da8fd9b0ec70e5d;
mem[18] = 144'h0819f8db0e71f67202e70e6b02ddff100d2e;
mem[19] = 144'hff71066d073401a50ccf0b66f7300b78f5ca;
mem[20] = 144'h0961040bf9a6f961fb32fd570604fe85f078;
mem[21] = 144'h0ea30e07fdecf329f9dc0d1e0f0b0396f57e;
mem[22] = 144'h068b00aa0edb0fbb0c1700950c5808a80bd3;
mem[23] = 144'hfa570f8afb38fc97f3d90041f1170f77fd65;
mem[24] = 144'hfa42fda3f666f711f3de0c8502d0f75afb68;
mem[25] = 144'hf26bf050035ff265fa0bf2ecfc91f7f00d7b;
mem[26] = 144'h0d8f0bbafcc5f139f8c9fdf20b1f0811f80a;
mem[27] = 144'hf3070a68f9a400fc0d440f0c042c081201ed;
mem[28] = 144'hf5c9f0970280feedf086074a061f0a51fffe;
mem[29] = 144'hf20107b3f3f6020208c60e74f5c505bc044f;
mem[30] = 144'h0cc6027308d00380f9140433f0ac0a9afc4b;
mem[31] = 144'h0412f888f70c0d9703c6090a062b06d9f921;
mem[32] = 144'h02d5fd2c005cf831f0110e05f5a9059bf9c7;
mem[33] = 144'h055afdc302350145fbcff132fa600b40fc10;
mem[34] = 144'h0bc80ecbeff3f4350033008509c6046bf023;
mem[35] = 144'hf1ae0823f543fbedf4fdf7300f650295fdf6;
mem[36] = 144'he9edef29fd0503bef6230575ff78ecb3f366;
mem[37] = 144'h03f0fa82f048fa190d8501fcee2d011bf141;
mem[38] = 144'hf0900801091cfc6dff63ff5105f4fd7f08e9;
mem[39] = 144'h0773f7d5e65bf2ccff4bfc25f9aa025dea2b;
mem[40] = 144'hf167ef7cf26b08dbf68f0578ef92e834f311;
mem[41] = 144'h0b26073d0a9d0155fd450887f77f0832f517;
mem[42] = 144'hfe3402b202daf3bff7b1f62cefe6fe7bfbb9;
mem[43] = 144'hf6bafa57ff53fe5cefdf0a700f170065f357;
mem[44] = 144'hfdacf4a407f4f6c7f824f9acf8470d96053f;
mem[45] = 144'h01b700190e94f62005de092ef134f242fb0a;
mem[46] = 144'h0647087ef02f0703096f0a5d057708370bb7;
mem[47] = 144'hffbc09ddfa35ee7204970887f68901a00671;
mem[48] = 144'h05d7f8590d14fc10f8ed03aaf241f0d4015b;
mem[49] = 144'hfc65fb3ff6dbf51a0ccfff1001e8fec3f049;
mem[50] = 144'h0b630c4befcc0a46f6f9069f0141fb7502f7;
mem[51] = 144'hfaa0f732faf9f5a50b6c0a78f26402aa0004;
mem[52] = 144'h0438f415f471f625eeb2035ef255f58601c9;
mem[53] = 144'hfd74f504093b0dbe086f0b6afea0f6af0a28;
mem[54] = 144'hf7060fa40b93f7aafac2fe70fd5dfbe90ac8;
mem[55] = 144'h082803ebe722f19ff8fe06e505c7f62007c3;
mem[56] = 144'h0274ea25ea88fa7204ba038d0ccff21bebc5;
mem[57] = 144'hed78ede10805feadfc3cf1b302fcf372ef9b;
mem[58] = 144'hf95a062807c4f90e0ae80b400a8c00540b57;
mem[59] = 144'hf29cf06f0765ff06f40df65708ab018704c1;
mem[60] = 144'hffaaf83df49c0dc80706f182fd6805e60953;
mem[61] = 144'hfc61002c06890a560bdffbfa01d003150d43;
mem[62] = 144'hf3a70e05fe85097f0c6df668fa1deffaf0a4;
mem[63] = 144'h051cef29f1b2efd8f437f487efe20beeeda7;
mem[64] = 144'hf35ff988f2e1fefffbd5f7fef4ac0193ef46;
mem[65] = 144'hf6fcf18ff71df9a2f9e1fc170a73fc1cf727;
mem[66] = 144'h0b43071cf03507580e6e098f09ddf247ff67;
mem[67] = 144'h00d10bd0f987fd500868fa4b09f3f12a0430;
mem[68] = 144'hf93aed80ffbe0a79f9f002cff544f34afc13;
mem[69] = 144'h00b8ed84f0440128f13ff761f2f9f1ee07b4;
mem[70] = 144'h0a4c044201650579088b076a09b10c330902;
mem[71] = 144'hfe90fa850921fd880b670360086c00bbf29a;
mem[72] = 144'h049d04e3e77afafff39cf32cf55ae5d5f33e;
mem[73] = 144'h00e9f653f563effdfc9bf1f2026301350c8b;
mem[74] = 144'hf73506d2fe6a054f02aef8c5ef6a01910018;
mem[75] = 144'hf26f0517077befa2061afbcbf260f8f10513;
mem[76] = 144'h0c7105a1f7620737fb160686fb94057b0748;
mem[77] = 144'h0e1900bfee88004d0001f480f150f285fd8f;
mem[78] = 144'hf9c6f9b50128f14104c9fd15065a0da8f060;
mem[79] = 144'hf6f5fe34fce005a201dc0990f85b033dfb77;
mem[80] = 144'hf307fe410c35f142f4adf3470a6c0ab6f5a8;
mem[81] = 144'hf7b2fe020a62f9090e390101fc87f3f2f0d6;
mem[82] = 144'h05b6067dff770c92fb97f663f124f3cd04fc;
mem[83] = 144'h02f7fa2409e7ff530408f00e055cfecb087b;
mem[84] = 144'h0654fdebf0b8fa69fb5cff2a02a3fec8f9d9;
mem[85] = 144'hfb40f84debb707c3f02df5550034fe33f3dc;
mem[86] = 144'hfee6f6120cdafbfb0e20ffd10af5005d0f25;
mem[87] = 144'hfcc2059ef590f0bbf611f697fa4503c1eec4;
mem[88] = 144'hfccef31b0265eea80b1ef63ef5b1f4d7016f;
mem[89] = 144'h0b8108def612f35eefe007c3f944f72b09fe;
mem[90] = 144'hfa6ffaffedf3046a01ad06310ee506360dfb;
mem[91] = 144'h01e6f77ef9e8f21d0999fdc106c108b9f71b;
mem[92] = 144'h0119ffbcf14ff16bfaec061f0bd1f6c5f4e3;
mem[93] = 144'h017a00780b7f0285fc33070efbd10cd8f6d1;
mem[94] = 144'h05eb024d02d704ed036b0eb5f017f4a1fa89;
mem[95] = 144'hfad4f5acfd6101710a340781f20d0c6e09fe;
mem[96] = 144'h031af78bf3f4f739f24f017af9a1fe4d0713;
mem[97] = 144'hfc400319fc720b01f0b00fc403df0d6d0b52;
mem[98] = 144'hfcfd04a30c1bf4e1feaaf36b0b250cf0fab8;
mem[99] = 144'h07a4f48d0daa01eb03b60690fbeaf33507a2;
mem[100] = 144'h0463f757edbaff0ef60f0cf80bac03e2f1a4;
mem[101] = 144'hf3dbff3f0a88f1900c31fd2a0baff7d3f8a6;
mem[102] = 144'hfb42f3caf2a002650457f4bdf570f64bfa0e;
mem[103] = 144'hf8650b4b0488ee56ffedf672fb93efddf0d3;
mem[104] = 144'hff40f7ea04aff7cf0b750dde0a70046ffbdf;
mem[105] = 144'hff4bf0ecf7b9f2000b1904ebfc9e0cae0881;
mem[106] = 144'h042bf16c0fdbf583f66cfab6fff6f87a0577;
mem[107] = 144'hf2a10b4206f901f509f90cfcf08dfdba026b;
mem[108] = 144'hffb6fed9f1a5fcc5ef5bfcd8fa9f0580046a;
mem[109] = 144'hfe6cf4d7050df4aa011df03a055f0925f380;
mem[110] = 144'hffe8f351ff8bf498f0faf20b0e9f0b4e05ad;
mem[111] = 144'hfd40f8db0f3efc69f8d6029b0573f5b9febe;
mem[112] = 144'h09bfefd2f53af3abfe97fdfdfc190430019b;
mem[113] = 144'hf0ebf955f22d0d42fcc70cb50ed2effafd8b;
mem[114] = 144'hf109f254fc7dfd7e0a9503cbf374fa9af04f;
mem[115] = 144'h03e8f522f760f78ffeb8f3820b3e043ff7e5;
mem[116] = 144'h02feefd0ebf9fee2eec308ed08a40a8dff8d;
mem[117] = 144'hf7a2f0ca0d39fd3dff8b0a89fceffb92f676;
mem[118] = 144'hfce6002af12b06c30deb051efa4cf843f721;
mem[119] = 144'hfd3904820ba106d5f10801f1075fed930b03;
mem[120] = 144'h0035fa950585089804fa0e36009af355fc33;
mem[121] = 144'h06d5048efbfefb29fce40bf7042506f101ae;
mem[122] = 144'hf311034f0941fd320a5a0499fc450ade077c;
mem[123] = 144'hfae90a72fc240d93fa1e0eadf73e0ae10e63;
mem[124] = 144'hfb6d0c3f060b061ef8b4f540f4e8f0450aa4;
mem[125] = 144'h0098096b075ef6b3f435ef5a0dbeeec704f8;
mem[126] = 144'h04d30aa5f8db0019f4defd21f21d0c610ed5;
mem[127] = 144'h07d30df3fd2feeb9f5de02b7f7b40d0ef5d9;
mem[128] = 144'h0a10051104aef326fbd4061c04d1f9aff665;
mem[129] = 144'hfb16fcfff62c03e30655f0640a81f5eef2ec;
mem[130] = 144'hf79f00e101f6041f094df0b6f4d3f519f924;
mem[131] = 144'h04faf4670f21012af4a8f08cfc350878f5af;
mem[132] = 144'h0ea6f83f0d7e022cf818f3eafbf5fd7503f3;
mem[133] = 144'h044bf58e06fef2050adcfb1bf54ef12bf595;
mem[134] = 144'h01e9f337065f06a3001709ce020df8dcf5f3;
mem[135] = 144'h06250c19f06cf5df0ef4009af3c908a604ee;
mem[136] = 144'h08340c70ff2e0316fd760e63f00cf1e1058d;
mem[137] = 144'h0177f87ffe320470f17a0443fb0c0092f3fd;
mem[138] = 144'h08e5f20b06a408f20354fe25fde80918fcea;
mem[139] = 144'h014f0f3600df0879fa4f0185070b05c6f6e4;
mem[140] = 144'hf60a03bbf36e021bf27c0c310d5f0493ff82;
mem[141] = 144'hf04608b9fef90de70853fb3afbc507b3fd7a;
mem[142] = 144'h0d0bf1dffcf4f276064908f306fc0d2e0980;
mem[143] = 144'h0cd105a206b4fe0d078df0cff197fdaafb45;
mem[144] = 144'hf2dbf513f40a0c680a5a08490a2603650ae6;
mem[145] = 144'h01a9f322fb410c66065008cc0a06fa3ef436;
mem[146] = 144'hf0610b3c0320030afe15f13307470bdf0dc6;
mem[147] = 144'h019d01c90271001602e501f9fda4f3280a19;
mem[148] = 144'h006409cbf0440bf8f255fd7cff5e0a00f3ec;
mem[149] = 144'hfdb604040695fd69f93ff2d3fb510d39f52e;
mem[150] = 144'hfe700a0ef3c80e110c5e0433f57ef260f000;
mem[151] = 144'h061af276f799f1da0332f04df3780a6f0ad8;
mem[152] = 144'h08cff26c0deaf92f0352fff20b28fbb30b1d;
mem[153] = 144'hf6f9f56209f3041c02090114f40b0990fdc5;
mem[154] = 144'hf8c7025c0473f34208a90759f9490e6afb1a;
mem[155] = 144'hfa4f09a8f53c0ef0f47efa940b9b005606fd;
mem[156] = 144'hfd3703b2ffa1f486fdbd0d57ef9af4b50f3d;
mem[157] = 144'hf94507bb0b620118fb550d0c0d5aef70efc0;
mem[158] = 144'hf7fef2e60b7e01e80d580187fe7c0cca0299;
mem[159] = 144'h047705a20de0f9760f140693f0caf6240afd;
mem[160] = 144'h076609a6f29af10f0131fcc80885f8ecfd8e;
mem[161] = 144'h01ddff360be90f620053ff870e90f195f7ad;
mem[162] = 144'hfc33f6b8f266f97503f8f3b1f67609b80998;
mem[163] = 144'hf9200461f5c1ff1cfbe0098f0be306e604b4;
mem[164] = 144'hf06807ed00cdfb54f840f98808e3f5fef643;
mem[165] = 144'h0bb00dad018c01310083086bf886f3c108eb;
mem[166] = 144'hf64a0a2904410851016dfe18fee5fc08f879;
mem[167] = 144'h0374f66bfef3f294fd8a04ab0425fa770caa;
mem[168] = 144'hf6baf9d70575f4220deb03e4effff81b0793;
mem[169] = 144'hfb5706acffde067ef2f50b3dfb2904aaf012;
mem[170] = 144'hf974f52b00e7fd3df55d004efa5109fcf9ae;
mem[171] = 144'h03dcf1930642f78ff9220c50f7bcf0c90e3b;
mem[172] = 144'hf7e402b7f6a808a9fa18f7d7001bfbb40465;
mem[173] = 144'hf81d05bdfaef0f14017701070cdd0b630232;
mem[174] = 144'h03c407a2fe77f662011d05e5f771f7a30708;
mem[175] = 144'hfae40baaf62308000653f4740f6df982f41e;
mem[176] = 144'h0cecfd1305140ad70a250228fbf909950165;
mem[177] = 144'hf223f95b0327049d037dfc74f5dcf4a0f717;
mem[178] = 144'h0d070a73fc8709060e930a32079d077efa8e;
mem[179] = 144'h08c8f7b7fe7c022afdbe05a20c4a05c30345;
mem[180] = 144'h0a7bfb6cf5a60e6df590f3e6f700fc5204c3;
mem[181] = 144'h05f00a7102fb0b22f61c0c7b0f4f00730533;
mem[182] = 144'h0adb089d0f09f5570a1df839f5d5073ef860;
mem[183] = 144'h07b403d5016b078b0c45f7cc093b04fef01a;
mem[184] = 144'hf4b80d08ff1dfbc7fe0df0440976fd190aeb;
mem[185] = 144'hfc16fbdf01090fb8f4a8faae08730cca0418;
mem[186] = 144'hfc9906d4fb6008caf34c06bc0f93004b09f5;
mem[187] = 144'hfe540c4ffa7efadbfcfd066ff43d06abf147;
mem[188] = 144'hfe0d0e88fac2f1860d2402f60b3604880970;
mem[189] = 144'h0a7ff3360194fa3cf37f0d63f84bfc7cf445;
mem[190] = 144'hf933fd2a07f7fa1d0c810199f3ed0deb0ea3;
mem[191] = 144'h0f2df7e4f533f04ef1c10d75f16af27006a3;
mem[192] = 144'hfe78fa76f0dcffeefeb7f690f613097000b7;
mem[193] = 144'h029bf061f823095207c50a26057407470b9e;
mem[194] = 144'hf9aef69afaf1fbe2053afc0f0bbfffba069e;
mem[195] = 144'h001b024ff2f2faa80184f860f66ef0c8fdc6;
mem[196] = 144'h03bc01b6f3b9fa54faf9f8d9f4d60143f98d;
mem[197] = 144'h022df950f18ffabbef7ff48b0bab07e1ff6a;
mem[198] = 144'h01d40813f9d4ff8d0b86028202c2fcde0cfb;
mem[199] = 144'hf2f1fb6f0421099e0acff79b05afff15fa2d;
mem[200] = 144'h0105f772f3baf9920f82fa7aee8ef49cfcf9;
mem[201] = 144'h05d2fa01f38ff1f0006803420b36093e0261;
mem[202] = 144'hfa18fbf20698fdaa0106fed20fd806f2001a;
mem[203] = 144'h06b2faa209e60af60dc70f5609bc0e2efc13;
mem[204] = 144'h0c7701f3f954ef3a00550322f73e0650f2f0;
mem[205] = 144'h09e6096b0556f08ffd4cf60902e4f05704b8;
mem[206] = 144'hf7630c4f032b0b97f2070b72fb220e4af87b;
mem[207] = 144'h013df07c03f504ea09640d4dfd92f70b09e7;
mem[208] = 144'hf1df078e0f17f2d4efff0e2e04320d32f3e5;
mem[209] = 144'hff080ae9f8cff99408730b790761fe4406bc;
mem[210] = 144'h0b5fff17f7cb0e9ff87cf755f664fc770174;
mem[211] = 144'hfcbff94004010a730a99fe3307460bf00185;
mem[212] = 144'h0229f6ec0150f2a7eb28f73cf62e07c6edcb;
mem[213] = 144'hfb3fef6504ba08430c4004c402b4f78affd7;
mem[214] = 144'hfa77061000e5f77808d5f95c0757f591fda0;
mem[215] = 144'hf8ae0123f408f042eee6051a076bf180f93d;
mem[216] = 144'hfe7b014501e40b250880efcffe84fddbe0c0;
mem[217] = 144'hf451ffb4030dfce807530332f07cfc08f3fc;
mem[218] = 144'hf640f6660e11faa90a56fe14f0990385f272;
mem[219] = 144'h025ef179f9d6f12bff9d0e0a04e5f6770699;
mem[220] = 144'hfa06073bf3520af8f81aef9afe84ef790b8f;
mem[221] = 144'hef4a02a70742f403f305f4c70083f5e6f43c;
mem[222] = 144'hfa21f3d6fa39f50ffd56fa1905ea0eaaf300;
mem[223] = 144'hf8ae0ac505abf1be080ef9310036f75ff2a6;
mem[224] = 144'hf7950637ff3afebdefe20065f016fe05f26d;
mem[225] = 144'h04fff5e30c0bff1cfa5b0fde0a27f944f99d;
mem[226] = 144'hf3c4f8daf357f56e0703fbc707460b96f043;
mem[227] = 144'hf2f0056206d40404f243f3f104a7ff24fa29;
mem[228] = 144'h0579f55a0053001ef28006c10eecef1df8e4;
mem[229] = 144'hfdf9f35d07d4f584ff74ffc7f9230339f6f4;
mem[230] = 144'hf2eaf7e2f9960b6a088e0a3c046e00880f26;
mem[231] = 144'hf3f7eeddf599fdbff59a0a62f826fefffa2e;
mem[232] = 144'h05cdf061f32a086afbf8ff7dfa9af0bff7e7;
mem[233] = 144'hf588fd39fed8ef660766f3c90a990a100bd6;
mem[234] = 144'hf6b70b860834f0f7011c0159fd590435fc89;
mem[235] = 144'h04dd0d83fb4501b7fa630a060875f3690ded;
mem[236] = 144'h0f45f8a4f4cef1aff0f101ab01170dcafb52;
mem[237] = 144'hfb66072cfef5fcd70ad9f3f70aa3026a06dc;
mem[238] = 144'h0111f988fc26090afa06f6bbf4980f8af598;
mem[239] = 144'h023cfa66ef8e065dfb5a016101e1fde90da6;
mem[240] = 144'h0769f501fb470307f53ff8b7f909fe83febe;
mem[241] = 144'h092005950c80f1e0019bf61c05c8f78bfc1d;
mem[242] = 144'hf9c8faa7f37808f301f3f595037df5a5fd84;
mem[243] = 144'h0a79f9fefe30f8890e4d00a60388f5cb0aa2;
mem[244] = 144'h00d7f741080e056bf708f523012cf1af0a70;
mem[245] = 144'hf8730381088ef0eef23e0aa30118f1aff95b;
mem[246] = 144'hfbc10991fa6f050b0bb5fa37f190f150f04c;
mem[247] = 144'h07dff474f16d09c901adfa1af136f8220aec;
mem[248] = 144'h0115ff05f336f6400c98fc8cf892fa71f7b3;
mem[249] = 144'h0bbf01f6f7d904e70c4d0db10819f253f49c;
mem[250] = 144'hfbbff2060b1bf2a00750f2aa012ef505f733;
mem[251] = 144'h0e560b16fc9705220e87ff1ef9a9f0a8f4e2;
mem[252] = 144'h08210a5cfb53fa82f0410212f357f475041b;
mem[253] = 144'hff6af0c10a4cf946ffebfb5cfdb1f3a3022b;
mem[254] = 144'h05f60bb00f7f075b0125fcbf09460a27fbc8;
mem[255] = 144'hf59ef9330b3c05290996f654fa75f2b6f39a;
mem[256] = 144'hf145f3b60679f2c9fba8f751046e0330f0f1;
mem[257] = 144'hf613f4bdfdf809710b190b8bfa8efe6402c8;
mem[258] = 144'hfd4f0da4f8840b0a0f2208ca00690d91f0e6;
mem[259] = 144'hf443fd9604330cae0a0ff589fc8c011ffdaf;
mem[260] = 144'hf1d4fd08fe39fe270057f1b505130c8cf86a;
mem[261] = 144'h0e0e009ff28a0c8afdbff8a607aef0010a1d;
mem[262] = 144'hf1d7fc8a03760563f087018005d4f2af0b0b;
mem[263] = 144'hfe57f86ef523f152f4690bbfed12f9a80a5a;
mem[264] = 144'hf75efa1b0597f1bdf5f2088effb8f96a032c;
mem[265] = 144'h032ffeb1f6900604f6adfd940577ef3a0234;
mem[266] = 144'hf233f3620fcdf2b9f468f046f9adf901fc82;
mem[267] = 144'hfaa309980eadff2809e602bc00cef3bffa60;
mem[268] = 144'h0ae1ef95f1a3078e064dfad2f729ef90f583;
mem[269] = 144'h0f00f0cd0948f996098af4860cc6fd59efbf;
mem[270] = 144'hfc2704690933fe20067c0a0c0830f78d0b94;
mem[271] = 144'h05240530fa0cfec70d48080a0c9cfe01f85b;
mem[272] = 144'hfd95f5910e510f4c06fa0e7e02f20af6fdea;
mem[273] = 144'h0ec40f2df89afb2e02ccf9d4f11cf5ef011c;
mem[274] = 144'hf6b9f0f6f883fec2f9a0fa8f0eb20a4d0915;
mem[275] = 144'h0887f72506f2f077fe1205e3f4ac060dfeb8;
mem[276] = 144'h01c6f11f09690690f3abf08d058906310841;
mem[277] = 144'hf28ff8f20d3d06a007eff9acf298f256f1d4;
mem[278] = 144'hf6240bc80b9cf3a70f5f0cfc0527fbfcff00;
mem[279] = 144'h08d7fa970c67f091f870f322f47209da0414;
mem[280] = 144'h00c2f07d01eafea4ff93089efe700c1e0b74;
mem[281] = 144'h0886f4080840f393fca8f7aff90b067c05c1;
mem[282] = 144'h099c0bf80cf5f59af4ab02f9f861fc9406f6;
mem[283] = 144'h0e46f879f66304db0e82f74302580ef702b8;
mem[284] = 144'h031d0b6402bbf264fb500cbdfac20375f3ce;
mem[285] = 144'hf35a0cf00c48f28c0e2c0dd2f6840937fbe7;
mem[286] = 144'h081708f6fdbd0ee8fb120475002dfbf5f883;
mem[287] = 144'h07d20a8505fffc99fe820456f5be04250a52;
mem[288] = 144'h013001c3f9b303adf4ce060cfa57ef8200e7;
mem[289] = 144'h00f8ffbb011b0a41ffb3fd11f3acf92cf9ed;
mem[290] = 144'h077e05220cf004b7ffd9fa1af585055a0f1a;
mem[291] = 144'hf051fcc5f5a0f6860982fbacefb2f725f73e;
mem[292] = 144'hf0e8e631fb600aa5ee4f020e02b504d5faec;
mem[293] = 144'hfbecf680f860034bfe42f50405d9091ff853;
mem[294] = 144'h0dcff45df63402db0ba4f1b0f0a00de1f4de;
mem[295] = 144'hf798f500023e0914f1e10756008101ad089c;
mem[296] = 144'hf036f335ff32ee7cfd30eee309e4f84afeca;
mem[297] = 144'hf22908d5edbd011ef38efc9d03fef1890a71;
mem[298] = 144'hf60903b5ff5302710d6d0820fa8505b4fc93;
mem[299] = 144'h07c30846f2e1f629fcecfe3c0961000bf9b0;
mem[300] = 144'hf2d10a9af584ff68f7a405200324ff6ff6e6;
mem[301] = 144'h0db1fd2bf3f30e0e0003002afe9909da0883;
mem[302] = 144'h0e8c01810afdf03ceff6fbf50d040cfb024e;
mem[303] = 144'h0e52fd0dfe7e061e04140147f74e09500a90;
mem[304] = 144'h0e6209a605b5fd5df8b806a00f9bf5b5040a;
mem[305] = 144'h0d090beff4c50f190ad709f6f8e5f7760a85;
mem[306] = 144'hf6d8fb2ff5e8090bf913072ff64ffed005ef;
mem[307] = 144'h06b7020af26908d5f84af63ff673fc6dff55;
mem[308] = 144'h0757f66efadc08e3fb84f5c1f15c055a0522;
mem[309] = 144'hf16000c3f89205c20c8ef317fdb908d00c93;
mem[310] = 144'h08ff0d9ffbb6fb460463058207ddf205044c;
mem[311] = 144'h00d6fe8dff56fb74faabea9f0535f275fda2;
mem[312] = 144'hf17b06c3f23905180087f3e3ee2eecc1ff7d;
mem[313] = 144'hfe65ef5cf3a00c00f4fc0955f04308bb0318;
mem[314] = 144'hf5bbf1ec0d86044604aef54c082402240366;
mem[315] = 144'h0cebf50905def5a5f3e401680b33026a0b6e;
mem[316] = 144'h0d31fef10cedfb220b9c0a6709b7fa00f3b3;
mem[317] = 144'hf7a2f9fef0c7ff70079effa1f0dffd36fb99;
mem[318] = 144'h0accfb42fac302cbf3dafadefafef0f1f361;
mem[319] = 144'hf39a02450804f2c6f8420cad05fd0620075c;
mem[320] = 144'hf692fcecff630963038e04ecf3dc0bc3efa9;
mem[321] = 144'h045f05f1095dfe950580fb7e0a8f08e9f75a;
mem[322] = 144'h0a2cff7affaff5f7f24b02b704690bf908d9;
mem[323] = 144'hf8b6f0cefcb2076efedd010bf2b5066ffeae;
mem[324] = 144'hee7ce90cee7ff32de94fee40fc94058500d2;
mem[325] = 144'h092505460b94ed28f9220b9ef2c7f7c3f13a;
mem[326] = 144'hf256f39ff5c1fcc606360619ef8e0bd7fae7;
mem[327] = 144'h05cafc75ee82028700a7064efe27effdf717;
mem[328] = 144'he81debd5ee2ee414fb05f54cf56500e1037a;
mem[329] = 144'hf5a2f730f0a30b01fb5908300db1076a0071;
mem[330] = 144'hf6c3fd6009dcf25d0b5af629f4a6efb6f610;
mem[331] = 144'hf6850073f09f0b99ff6f03d706020634014d;
mem[332] = 144'hf88a0586098b085606b90a9dfd300b84f3bb;
mem[333] = 144'hfae6f647ff20f5a90a45fa3005a20aeefd56;
mem[334] = 144'h09f5ffd4f2bdfc71fedbf71a086bf65dfaad;
mem[335] = 144'hede7f9890c30fb18ef4f091eef75f2ae0292;
mem[336] = 144'hf374f46307adf714f8d708da07600dcc05b0;
mem[337] = 144'hf4deffabf639fa8df2fdfd370cb305c20cfc;
mem[338] = 144'hf91cfa3af3fc0790f37508e307770e81025f;
mem[339] = 144'hfce3f37f0e88f83f05def264f6cc0c6ef32e;
mem[340] = 144'h0d390382fe610c1afa9006cefa26f7c60a1a;
mem[341] = 144'h0a8804d2f0800107f34304adf189052a05ce;
mem[342] = 144'h0de2f061fdc4f55e0d480db80bbbff16f286;
mem[343] = 144'h05d3f2aaf20909e3fa0707ebf151f47ff14d;
mem[344] = 144'h03a4fbb9fe2ef2e305e80166f3d2004ff6fb;
mem[345] = 144'hf9b7f5e40242fd97f6dcf83e0a3c02f5ed92;
mem[346] = 144'hf13f05a600b2051d00240c38eed9efc0eff4;
mem[347] = 144'h03950a080270efc4fa4d009af15b00100eba;
mem[348] = 144'hf8e007d7f47d0a360ce9ff64efc70e0cfe66;
mem[349] = 144'h0405f2e30569f5dbfab900520813f5ddfa43;
mem[350] = 144'h0bc8fdce05cf0e42fc2b076e0398f9c6f1d7;
mem[351] = 144'hf5590e0507b5f4920e2a04c2f0cfef7301f7;
mem[352] = 144'h048e054300fe09bcfa4b0293f4c0fd11f47a;
mem[353] = 144'hf19c0340f4e5f118000ef2ebfe39fa32fbd6;
mem[354] = 144'hf5740ac70d170d6ef268fb81fbaff0b7f91a;
mem[355] = 144'hf126f39c0ace0986fb1ff88d0dd5fb5f05cb;
mem[356] = 144'hfa03fa31f834f3840a6a007c006bf673ec83;
mem[357] = 144'hf5c6f1ec0564fec109d6091f0b65091df077;
mem[358] = 144'h034bfc53ffba0a83fdcf0ea1063df7c8fb3c;
mem[359] = 144'h057d08e5ec82f1b3ee43035cfcbf0489f09b;
mem[360] = 144'hfc7cf786e80903f6f863f8daedaee479e6cd;
mem[361] = 144'h0bd90b75f8870f8a02000c0f0930fcc9084f;
mem[362] = 144'h06d8fd2f00410f23fcea017dfdf7f1cd01bd;
mem[363] = 144'h0bc1f5f3f696f75cf1ac016ff9080e56f76c;
mem[364] = 144'hfd9df16904a3009dfc89f252f5a0f22dfe83;
mem[365] = 144'hf52a088befe504e9f1d6feaaf53ff4360d4b;
mem[366] = 144'h057300eaf064f75cf5a7f09d05aa095104f0;
mem[367] = 144'hf2bbf48ef21c05870829f21e05cbf976f8dd;
mem[368] = 144'hf3740cf7fc00fa7df4ec0019fdde09de02ec;
mem[369] = 144'hf075fb22f0cf0d25f07105510f9d027c05c0;
mem[370] = 144'h07290b550db10fd40fe0f5e90f3a0a4c07d7;
mem[371] = 144'hf962f2b7f0d00d67f7f5f249036ffc4cf60a;
mem[372] = 144'h0fd0f2060195f7090bc808e2037af8090b59;
mem[373] = 144'hfef9f6ccfb8501ebf4cf00d1fe31f19d0ded;
mem[374] = 144'h0590f91b08340dfb0cff09fff2b6f9670507;
mem[375] = 144'hfa2f00160877f409fa3f0bfd0a0d0b3def63;
mem[376] = 144'h009bf64a050908c4f14af648f63ef8430916;
mem[377] = 144'h0258ff2904560abd007b03b803fa0e0dfc66;
mem[378] = 144'hf6f80ce200b5f4c60a6a09c8f8d30beff191;
mem[379] = 144'h0df10f6500a5089708410116fac2fc100b22;
mem[380] = 144'h0c15f54c0ddef108f29507ef0534f0270720;
mem[381] = 144'hf35a09bffe460446fafef1800764f3760680;
mem[382] = 144'hf2e504c2049cfdf40a4ff38d01e3fa700233;
mem[383] = 144'h0298048bfa2bf7ab039cff4af73909ac0d7e;
mem[384] = 144'h0f70f6ef0b320e1ffc640c1d0a9b0daf036b;
mem[385] = 144'hf64000c8fa390658fdff0740f112f92cf8bf;
mem[386] = 144'h0e9a0187f45d0c41032f025bf11f05190633;
mem[387] = 144'h07b605300db90730f7d0fbf3035804e3f873;
mem[388] = 144'h0821fc050a8e007c0c2cff05f9a5ff960a73;
mem[389] = 144'h03eaf675f256020a0acf09c40bed0498042c;
mem[390] = 144'hf788fa6ef47d0c6c0f180b5efa8e02f9f448;
mem[391] = 144'h0c92f8ddf8bd0ad40033fa09faeb0dfafe52;
mem[392] = 144'hf5e90431f02905e4fb2903bff37800d3facf;
mem[393] = 144'hf457faf1f525fc22fa68ffaa04fbfee2fdd5;
mem[394] = 144'h03baf2bc068ef2e0f933fed8fd3df71ffdac;
mem[395] = 144'hfcd40a6007a5fe05ff71f841f6a901c7fcc6;
mem[396] = 144'h01e2ff03f200f775fc3e018a05880cee021c;
mem[397] = 144'h0e04f606f7740f96076cf9f6f95a032602db;
mem[398] = 144'hf0db0d9cfb590d560a41f847f8360611ff7e;
mem[399] = 144'hf7d2f166fdfc09820c85f77cfc8c0ea70b11;
mem[400] = 144'hf7eb091ff36ff6f70c88fc84fb6103a7078d;
mem[401] = 144'h00d108ee00fcfd720c8bf9710b64f77cefff;
mem[402] = 144'h0ba3ee5c0af80019093fff75f9edfdc3fe00;
mem[403] = 144'h0ca1ffba09a7fc3900660b23f6800beb031f;
mem[404] = 144'hf17defe1fc92f1def229fa550962ebf0f4fb;
mem[405] = 144'hfb8ff3510b7af5730828f66afb0b0847f1ac;
mem[406] = 144'h0d8b04660b7602b6fd8ef52cf383f2f80670;
mem[407] = 144'hecf6f7a6fd47f6d20c4e0670fd33f5c2fc88;
mem[408] = 144'hf90af79df2a9f14b04befbeaf687016301a4;
mem[409] = 144'hfb950c3df7e70bbdf630f188fbaf075af5ec;
mem[410] = 144'hf145f533edf6f708f4ecf1670b7e0b1ffd0a;
mem[411] = 144'hf1a500cefbd30074f515f53f0844f287fa99;
mem[412] = 144'hf8d40a1c010bf35af1c3ff63f3bdf7b4f993;
mem[413] = 144'h09060b4009820280fbe2fa93f907f9bb0a5e;
mem[414] = 144'h099cefd1fa4a0881f4c503810eb0fe79f6c0;
mem[415] = 144'hf173f623023cf8eef208ffeb0b31fc8a0774;
mem[416] = 144'h023af22303f70d010c0af7a6f1ddf852ef90;
mem[417] = 144'hf434f6fb08bd0d31f0b0fa9d0054f6760ca6;
mem[418] = 144'h03d1fc32ef54f01c0b8dfd7d03d40137fd29;
mem[419] = 144'h06f8073df3f5fdd2fc8e022506930989f290;
mem[420] = 144'hfdb8ff91e584f0d6009df652f3c80589f13c;
mem[421] = 144'hf04d06fb01ca089bfc440468ff0ff047faed;
mem[422] = 144'h00affb920e19fcc4f792fa40f59ff173fe64;
mem[423] = 144'hefa60263f96af24bea32fc99f9cdee44f11f;
mem[424] = 144'hf060e887f80b00420931ff4bfed6ff49fc72;
mem[425] = 144'hf702fdcbf0480243f959007507bbfd45087e;
mem[426] = 144'h063afd14edd4f254fe02018dee940622ff96;
mem[427] = 144'h09490980063f07fbfa52075a06a302fe0132;
mem[428] = 144'hefad0d3ef2db01f9fd5f0cef0030f964fc3f;
mem[429] = 144'h0abefa0bf7ebfaea0747fe340986024c05b7;
mem[430] = 144'hff91fcfefd30fe3a0548f2090e690e4a0160;
mem[431] = 144'h0050f7d6f6a80aa20b520667ee5cf805ede9;
mem[432] = 144'h0a1c0a9a0fe20043fc94f90101d1fceb0b57;
mem[433] = 144'hf254f93c099d06e10e0d07760f36059200ee;
mem[434] = 144'h09f90a630719f07b0a77fa27f13c0988f4cf;
mem[435] = 144'hf48ffc930f0c0b96fe10fb93f040fb9bfd34;
mem[436] = 144'h0b960bbf0c3ff7b6effff14bf01afa5cfef3;
mem[437] = 144'h064607590a59fa0808a10b17f29df2d90200;
mem[438] = 144'hf02b07d80e20f020040c08a70eecf38ffedc;
mem[439] = 144'h009ff033f1960a7603f00f34fc7dfb2407ea;
mem[440] = 144'hfed10487fb1e00420859f00df680f739eff0;
mem[441] = 144'hfadfffe50ca5f152f236f39c0358fcf50d09;
mem[442] = 144'hf0720edc07b1068e037304150b350780f284;
mem[443] = 144'h0d75fbc6f881049609a004c4fe02fb9ffb78;
mem[444] = 144'h0b640d6b0fc101eb0676076bf2ac03f1f126;
mem[445] = 144'hf277f237f1a90d54f03002b7f630f0d0ffb7;
mem[446] = 144'h0ec507d5f7dd0de3f2f5f223f7600954f0b4;
mem[447] = 144'h06f3fe58f27b06940b280eeaf76f0014effa;
mem[448] = 144'h09f00958f74a00fe056f0cd5f866fd17fb73;
mem[449] = 144'h0180fa58eff803f0f51e0f620bfb001b04bc;
mem[450] = 144'h0abe00de0b09f30b0dfb0f1ff43103b800c7;
mem[451] = 144'hfa1e0185f6fc0dc20dd703f7f25b0058f50b;
mem[452] = 144'h0366096ef6fef75206ac049af59df3edf488;
mem[453] = 144'h07a0fe060c88fcda0a18f15107ea020302e9;
mem[454] = 144'h0e490773fb8ff040029df0b20d91f06901b1;
mem[455] = 144'hfac5f034033afc19013af494eea0f80b03be;
mem[456] = 144'h0519ff470662eefcf829fdbefcce0bc4f63d;
mem[457] = 144'h06a4fd92f023fc94fd1c08f80a07f1e604be;
mem[458] = 144'hf2940565fb090edaf04f026efa07f10d0966;
mem[459] = 144'h0107fd85f3e306cdf51e0907f35f064f04a6;
mem[460] = 144'h0cfc07d10e85fb660e9bfc3ffed8070bf7fa;
mem[461] = 144'h0293f04eefa10d51ef8f0ae90dcd01aafaf5;
mem[462] = 144'hfa6c09be0a66f8f1f087fdfe0029f6eb0d93;
mem[463] = 144'h020ff30f0976089802a4f140f1f706210a8f;
mem[464] = 144'hffa30075066b0f31f7f4067af4350586fc8a;
mem[465] = 144'h0f500b5dfb96ffdafb260641f525f22502c1;
mem[466] = 144'h0c5af6e6fc560929f125f843f79f093cf643;
mem[467] = 144'h0c0df7d0026f015707b902ea0457088df2f1;
mem[468] = 144'hf207f565ff71f271ee6eeecc010af7c70aeb;
mem[469] = 144'h0555fdda02def52ffc000e56f38103aaf785;
mem[470] = 144'h0bdffa1508b8002ceff8f1140999f11a03a2;
mem[471] = 144'hee9cf65feddaff2b0798f7320504f32cf782;
mem[472] = 144'hefe7ff87075f0bb7fb37faa5f8b9f9c9f558;
mem[473] = 144'h040604eff27b09ed03b400aaeffafbca0f29;
mem[474] = 144'h018905760432fc840ca8f95400a6fc71f87e;
mem[475] = 144'h0ac4069ef5f80514027ef632064c06b6f9e6;
mem[476] = 144'h01f3fbe80a9df810079f0cb2fb9602e6f8f4;
mem[477] = 144'hf117efecf49603f60204f9e40d2008650b29;
mem[478] = 144'h0cb7fd6007a7f6d3087e0fe3ffcc0b17f22b;
mem[479] = 144'h055f09fd0723f311072e0b1b08980c4ef20f;
mem[480] = 144'h0857ff43053808a90e5d0b4c0663fee0fa64;
mem[481] = 144'hf536f2f4ffab0c02f663f2bbfb4ef1c507f9;
mem[482] = 144'hf75cfa58f7e101b5f47802250b7ff1e707f6;
mem[483] = 144'hf42e02e100010225f62efa3c0cc00c8809b6;
mem[484] = 144'h0d74fdb80304f4c90793fcf9fae40e06f9a3;
mem[485] = 144'h05d2f064f06df7fa0170060bf31ef1a00705;
mem[486] = 144'h045608140a77fef800e40faa0d73088ef83f;
mem[487] = 144'hefb70c04060a0ea7fe680ad9f7140981fe5e;
mem[488] = 144'h040bf2baf3470c750780f3e70ca1f1170a54;
mem[489] = 144'hf690f6f2ffe1fa41f5aa07ce04710345f4e2;
mem[490] = 144'hf653f79cfce5fe04f36ff79d0a44092eff93;
mem[491] = 144'hf92af4abf8e1fcedf0e4fc910f25f1bcf42a;
mem[492] = 144'hfa61f4e9fdc1ff09fb9d032f05c50943f18c;
mem[493] = 144'hfe17f16d0dfc06a3fbb5035bf4eafd6a07f0;
mem[494] = 144'hf10a07dff87aff120e7bfe4600cb0b31089d;
mem[495] = 144'h00400daef0a403d4fbcbf37407b9f1c70776;
mem[496] = 144'h0d480c6dfd41fa0803fcfc1dff890e7201bd;
mem[497] = 144'hf501f69cfee3f1ecf30eff0ff1dbf8460f65;
mem[498] = 144'h040af214f39207060736fb440d43fc7606e6;
mem[499] = 144'h0b3c0d2affc50c310e54f54cfc4f0d82fa6f;
mem[500] = 144'hf11bf07a0a1df88afa8e0c2df50303f4f31d;
mem[501] = 144'hfa88fd84ffd5f2530087f26002010e83fbf4;
mem[502] = 144'hf2d9f8970864f066009cf70a05d20734ffd9;
mem[503] = 144'hf0f3ff92fe7bf381f458f9e7f14cfb39fcc0;
mem[504] = 144'h089c0f07f1b7f39df72fff530adb03f4ffea;
mem[505] = 144'h0f0002d7f526fee00eab06d40edd033507a0;
mem[506] = 144'h057ffda20fec0a0ffe57fef20e110120f33f;
mem[507] = 144'h0ec1013ef3baf3befcaaf756fa510c960c3e;
mem[508] = 144'hf7b8f9feff340282f61601bc078e0f9cff26;
mem[509] = 144'h0b0ff7f7fffb09190aaa092c06470a71f9e9;
mem[510] = 144'h057a049400c3057efe0ff60c0b790aa90f62;
mem[511] = 144'h04920216084df76ff17b04cffb3dfbf00658;
mem[512] = 144'h0ccff212ffe3f1cef69c043ef5d7fb55f96e;
mem[513] = 144'hf53bf99bf146fea3fd85043cfe35fe0a0739;
mem[514] = 144'hf7cefbde0b0ff74e0be8f9fcf035fd640671;
mem[515] = 144'hff0d01e6f71a07dcf0d80d7d0886fd26fe80;
mem[516] = 144'h0fa20854008efa17f1cfeefb0382f8b0fd80;
mem[517] = 144'h04c2f78ff512073bf8c20d3d0e3ff2d907cb;
mem[518] = 144'h046af5dbfc1cfe580d33052204880c8a0b43;
mem[519] = 144'hf8bd0a8b03bb01b5f5e6f361f793fa0af824;
mem[520] = 144'h0e32f211f5fefcf70cfbfdc0f1930968fb1d;
mem[521] = 144'hf4e6ffd4f5df0e74fd7df34cf0ac0b55f45e;
mem[522] = 144'hf7fd027efd340e43f4f5fcc1f49a0c7dfba0;
mem[523] = 144'hfa0101daf1b4f9bbfb090f1b09540d9ef336;
mem[524] = 144'hf466f39afd2bfc2afc55f151faa1f32df8b7;
mem[525] = 144'hf5e600180a3af825ff440be9f920fab604f7;
mem[526] = 144'hfea10daf061b0eeefb10f39105e0028d07e1;
mem[527] = 144'h0407f88203eaf199f92cfca90cf006c1f60e;
mem[528] = 144'hf697fde60b13efd0f333f0d1f302f85df919;
mem[529] = 144'hf26efa520278f832f762008bfe00f8940ac9;
mem[530] = 144'hfd4bf5f10176f026fbeff04cf71002ba059c;
mem[531] = 144'h0d240e4af11eff76ef4affb20bd8f504f047;
mem[532] = 144'h0275f30ee7b8f2650577f87ff676f458fb90;
mem[533] = 144'h07f9f6d1fe92fae10a2f0c34fb50ec4d0496;
mem[534] = 144'hf1e6f073fa0cf025f498fe3aff69f5830558;
mem[535] = 144'h09cdf35803e4efa507bafa71f130f37ef9af;
mem[536] = 144'he74ae18ee663fbdbe990ff7ff6c9f32afa29;
mem[537] = 144'hfac3fe8dff93f3b00ab70207f1d20688f555;
mem[538] = 144'hfb48faadef700a7b09ee0d050cbcec4af452;
mem[539] = 144'hf4d00047069af3ecf29c0f30f2b60b1b088b;
mem[540] = 144'h042100200c37fbcc033e09900e7af5c8fe48;
mem[541] = 144'hf0d909f2fcd2fddb0d87f9390efbf12000bb;
mem[542] = 144'h03860a6ff8e80583f2dff8b0fd8b00d7f9c9;
mem[543] = 144'hefb8f896014c0ad1fa8ff4610d7cfadd0494;
mem[544] = 144'h010d01900c7a094701120d69f6390bbefa3e;
mem[545] = 144'h068206260105f451f27bf42cfa5d04460e12;
mem[546] = 144'h0849f71308c9f30bf69505610369043304e6;
mem[547] = 144'hff76ef66f3c20054f5bc0cf3f02af45df115;
mem[548] = 144'h0a31006108e6ef2c063e03d9f8ccfaaeee37;
mem[549] = 144'h0b07f2a3f9c20191fab7fb6ffeb003100d47;
mem[550] = 144'hf86bfc650e5c073302cff8590db2f87b0018;
mem[551] = 144'hf7a2075aec650a080aeaff660194f0ea0496;
mem[552] = 144'h0aa5ec7ffbe6f8d1038d01ef0bca07c4f24b;
mem[553] = 144'hfc98fd78ee96edf602c8ff0e025ff84ef6c0;
mem[554] = 144'h0161f89100b5f78f02c3f0ce0950fac5fe45;
mem[555] = 144'hf5600eaa0fa205dff2450f8e03e5f4cf02ec;
mem[556] = 144'hf5e0f957efccf19df15ff059f53902a5f400;
mem[557] = 144'h07e70274071c0728fb96f0a2f3d9fd960ad4;
mem[558] = 144'h044d00ce0bc60c240379f021fd5ef1b20765;
mem[559] = 144'h051e023203fa086109aa08130690fa45fb5c;
mem[560] = 144'h08e706b8072bfb85f7e4ff00f425003b02d6;
mem[561] = 144'hfdea0b48f6def182febef8a30d1a0cfd06be;
mem[562] = 144'h0661fecafb77036202670c570f410c230c37;
mem[563] = 144'hfe53fc8d02ee02a1f860fd5bf9b7ef52f82c;
mem[564] = 144'hf11109f60aa907d5eed30229fb850065f134;
mem[565] = 144'h06ea056c0291f0db0bab0187078307d7edec;
mem[566] = 144'h025e05480761fbfbef68f900062df6d507e8;
mem[567] = 144'hfb91fd9af48706caf167eb92ef10f3bcf98d;
mem[568] = 144'h057707db0498ee1b01baf2fce870e602eb51;
mem[569] = 144'hf00902cc047002020f14eed2f5b70179ef04;
mem[570] = 144'hf54c0958fb1c08ccfaad076f00e1eed1fcc3;
mem[571] = 144'hf380f618f7a20537ffc704450cc9f98d0d07;
mem[572] = 144'hfb410e30f2590151f0c8fce6f684f7e10703;
mem[573] = 144'hf7d1fbcaf3ab0a34ffb3f728fad2f13d07ab;
mem[574] = 144'h04edf73d09cd01ecfbc1f7f80d5d0ae0faf7;
mem[575] = 144'hf883fac5023507d4f4a20ac2f765f3d8fc86;
mem[576] = 144'hf617f740fc27fc23f21e00a2fa1107320476;
mem[577] = 144'h003af18ffd420bf1f7680f67ffbb0857f416;
mem[578] = 144'hf7c2f2f4f5d7f074f0d2fd7b0f460374ff9e;
mem[579] = 144'h0adfff7005d0f94ffb5e0cce0e510edff986;
mem[580] = 144'h0596fb400978f3b20d2ff474ffe8f829ff78;
mem[581] = 144'hfe72f9600a47faeefef309e00208fd32f8f1;
mem[582] = 144'hf0af06cbf17f0d8009950d97fba4efebf2dd;
mem[583] = 144'h0403fdbdef0d004cfaa5ee82fbedfe6d0144;
mem[584] = 144'hf711ffca0db307e2fefdf7160c5cf586fc8c;
mem[585] = 144'h0dc5051efd5d0ad60b78f76d06f804c8fc04;
mem[586] = 144'h00cd0a52f9430f5ff92d04f6f969055efdf9;
mem[587] = 144'h0c9ef62b0cbdf082f933090df1fffd330a20;
mem[588] = 144'h062f0924f5e5f972f02a0a330906fc930f21;
mem[589] = 144'h073a01e6f3b2f0ad0612f3bf0975fca2f93d;
mem[590] = 144'hf351f80d05b1fedcf199f2f2f1520ef30af5;
mem[591] = 144'h0727fbf20e57f10bfa3ef86c037f039e0a70;
mem[592] = 144'h07cef017f0b50076f4fc08770e53f3900f78;
mem[593] = 144'h034ff232f3def200fad1090506b40423fa04;
mem[594] = 144'h075ef1d0f0220deaf1630b7903b5038dfadb;
mem[595] = 144'hf52906350ab1fa060a8f089b012a0cbdfa14;
mem[596] = 144'h0a720488fb48082af9e00ebdefd3f978f61e;
mem[597] = 144'h086f03fa0719f3a2fc8bf1c0fe200ae0eef5;
mem[598] = 144'hf46bff2204f801e902540b3df1cef2f2fe84;
mem[599] = 144'hf89d019d06d8f882f8aa0492020f0778f8cd;
mem[600] = 144'h0d390149f9470c3def6df3e20a9f09a9fb80;
mem[601] = 144'h092a0b3ef2f402e0f825006bf7ebf20af00d;
mem[602] = 144'hf49c0ce2074c06d3ffd205ce07920b3c0e09;
mem[603] = 144'hf4ecf59bf16f0ba603ccf0e4fc6efc41efc4;
mem[604] = 144'h0192038d0c27f3540a90fa2cfae302440369;
mem[605] = 144'hf2ca0f6ffb6e094702220f14f9fc0d2cfe02;
mem[606] = 144'h0df6f0bcf35ff7d1ffd408f80bc8f1d207ec;
mem[607] = 144'hfbaffe100ad9f6190148f1dff7b3f9a2f74a;
mem[608] = 144'hff37f46e02a20c8cf195fac20107fe7e0e38;
mem[609] = 144'h0c42f072f9960eaa01c90ddc0544081df0ea;
mem[610] = 144'h0d0c0a1df2bf0ffc0dde0e550e570c0d0ecd;
mem[611] = 144'hf8ce0610f896f4b60e1affcc0b2f08d204e9;
mem[612] = 144'hf757fe56ffcd0e26035a0c10f3c3089dfcf8;
mem[613] = 144'hf8c3051dfbf3fb5a06550b9bff1f0a1cffc3;
mem[614] = 144'h074ff42d096a0beef90cf321077104b707c4;
mem[615] = 144'hf5e4fae4f0160cc40867f1440005f6cafcbd;
mem[616] = 144'h0072f02afbe40116f24a0110f951023df825;
mem[617] = 144'hf84bfce60db8f740f98cf82bfcc3028efb08;
mem[618] = 144'hfeafffe7fb47f690ff6af1680b990ec108c6;
mem[619] = 144'hfbbffb9d08b304d0f59ffa2f0b0ef334051c;
mem[620] = 144'h038df05ef3250f0cf5cef613f550f5d7f3cd;
mem[621] = 144'hf578f34503daf0e500540523fbfcfc51f845;
mem[622] = 144'h0fe209e9fde7f8b209160e9cfa70f579fd6c;
mem[623] = 144'hfd4605bd0b88fafefa010ad4f554fa7af635;
mem[624] = 144'h02950825018dfcf705b60404f7e2f227fb14;
mem[625] = 144'hf3d7f5f5080e05d50122fada0a9807ba05e2;
mem[626] = 144'h0acaf1a2fa74fc17fcdafc09fbe5086ff3ec;
mem[627] = 144'hf4590e9fef6d0607f122efd10a8e0809fc4f;
mem[628] = 144'hf38afd360370f9880153059af41e0440feb4;
mem[629] = 144'hf1630028050efec109f1f4f6f9fff49c0df6;
mem[630] = 144'h005704ff06cd01aef712f3f7ffcbfa620bec;
mem[631] = 144'hec8ffb1907b1fc8503bef6910aa3ec68f1ff;
mem[632] = 144'hf72e005c0de0087efe36f10befbf071c05cf;
mem[633] = 144'h0b78021f01cb0e3c0730fd19fd8dfe7eff7a;
mem[634] = 144'hf7c3053cf2e806850b22f777fe42f92bf4a3;
mem[635] = 144'h0787feb107920e8afbabf2c3feb1f7fcf598;
mem[636] = 144'hfaf8fbfbf4440958fa2d0a70fe730b0cf98d;
mem[637] = 144'hefd5f6da071d00d20dad0718febff0950f6b;
mem[638] = 144'h04a00584047e016efaae0617f33906c0f157;
mem[639] = 144'hf88ff6040f66f93b076e031d0028f3290629;
mem[640] = 144'hf8560f03fb5c033508e1fa75fdfb0527f611;
mem[641] = 144'hf946f0adf0fcf042fd4ff693f83c02920e79;
mem[642] = 144'h0f07f973f99e0c9e091cf681f74507f8f6ab;
mem[643] = 144'h08d8f83f0144fb48fc85f743071401340a1a;
mem[644] = 144'hf196f7600547f0eb0ea1f28b084cefed02e3;
mem[645] = 144'h0f1d01f8f13b01b5f5c10a6b03b1f349f071;
mem[646] = 144'hf61ff82bffbdfeeef2e3055f00970b03f2c4;
mem[647] = 144'h0391f91af17b07f5f7b0f8ac04de01620657;
mem[648] = 144'hf6d90011fe8ff369025af8200f8807f20eec;
mem[649] = 144'h04c6f786f87c03c605c4ff73efd0f6bb00d3;
mem[650] = 144'hf88ff75efa58f541f9c90c12ff19f0780102;
mem[651] = 144'hf9a902d903b2f68a0a2703320d92fbcc0bce;
mem[652] = 144'hf27b0794fa5e094b0d88f199fec00f040a36;
mem[653] = 144'h0f7709b9f147f9f6047af6b8f00a04bdf323;
mem[654] = 144'hfdd4f930f834f0cff87af387085901e7f69b;
mem[655] = 144'hfb99fa7a0c3d02fa0e3c00b7f967f7d109ba;
mem[656] = 144'hf2b0fa7c091ff22c09b4f9e2055904da0c0e;
mem[657] = 144'hf1f9fe6ff763ef3cfbd805af089608460699;
mem[658] = 144'hf4120754fe8f02e1f7c2f5bb01b9f289f48d;
mem[659] = 144'h0309009ff4d0028e0d20fdd40da6058309b8;
mem[660] = 144'h02a0ef83033f09450cff0a31f5a3ee760696;
mem[661] = 144'hfd5804d90510008209f20931f2a8fb7afdf1;
mem[662] = 144'h0ce2fb14073d02b9007dfcfc099afee9f938;
mem[663] = 144'hf0c5ece0f15ef54303bc090e0625f02dfc3c;
mem[664] = 144'hf97d0069f4aef806fb40fc2eff40ea140808;
mem[665] = 144'hf305fea0ef08f5f8f29b0292041e0b93fb83;
mem[666] = 144'h01d0ed7b05eaf8f60ec7f754efe8edb8061c;
mem[667] = 144'hfeb40cc10427f71c00cafd1a060c0f81f94e;
mem[668] = 144'h0d48fecffdbaf123f7a0fad4f4440e460dfe;
mem[669] = 144'h0c5a06830c3ff7daf5a000300320fe84fb38;
mem[670] = 144'hf10100080a49f68bf04f0c86f6ab07570ad3;
mem[671] = 144'h047f048a03650dce0e0af73cfebc0b690511;
mem[672] = 144'hf9850f950351faabf87604ac01820d18f8df;
mem[673] = 144'hf493f7b50f4c0aebfbfbfb49fd23fc630725;
mem[674] = 144'h0b68fe2efc530ab70379f9cd01e5f63e09ce;
mem[675] = 144'h040cf1560c21ef23f6460c00060ff13000a7;
mem[676] = 144'hf25103c10b0b0748fd660c54fff1f6e30b3c;
mem[677] = 144'hf4470cf7064808f202f7ffcc015c0ceffc9a;
mem[678] = 144'hf6c00ea001a20d7df43000300a6ef4acf3be;
mem[679] = 144'hfe22f4b7efb3f69808340376fbd4f15dfa0f;
mem[680] = 144'h0e3dfeb9f3edf67705aef5b0f81302ce03bd;
mem[681] = 144'h077009e5faa1058bf783f9f900abefcaf45c;
mem[682] = 144'h0791f72ff310f62300fc0a7e0b3ff30ff27c;
mem[683] = 144'hf1a8f28107280360f7c705b3f631fd71f2ee;
mem[684] = 144'h0a2b075305a8fe4b090300b4f99aefa6f3e0;
mem[685] = 144'hfb55f13706b901a70a12f8ac0aee087605de;
mem[686] = 144'h0fd70b1e008a0d19f3510eca0807f1350c58;
mem[687] = 144'h0dbe0cb802c0f7330f56f84af2d8f7d9fb44;
mem[688] = 144'h0d59fa7103f7f4a20cabfde0037d051f01a0;
mem[689] = 144'hf22c0d6ffe4dfef4f8fafe07f1c7035df594;
mem[690] = 144'h08620d200dfeff6f0c940b35f8fef3b8f227;
mem[691] = 144'h0766f80bf8c6f46ef17e0d38f225f1f8fad1;
mem[692] = 144'h08a6f059f753f7f2fc020ceef777f82aff45;
mem[693] = 144'hfbec0ecaf11d0a24fe2400a20d5d04bd0a74;
mem[694] = 144'hfb4af01b08c1f064088bf0270e4bfa58fffd;
mem[695] = 144'hf7e0030707d4f1e4fcd5f3060a1a02ee0005;
mem[696] = 144'hf41f0826f1dc076106370c5f021905bc0232;
mem[697] = 144'hf595f1d009fef4dbf03efdf30dacfce00b49;
mem[698] = 144'hfbfbfc9bfa77f2b6ffcafcb7fee8f782f3da;
mem[699] = 144'hf5330a02f6f9fcb9f706fb330154f89ef2d4;
mem[700] = 144'h0d8608affc6605140548f6aef1830c5afa19;
mem[701] = 144'h044508660f03f7c5fb9e0a46fceafb20f779;
mem[702] = 144'hf5d0ff680ffa0cee04d8fcaff32f0d230cf3;
mem[703] = 144'hf17305f60d4afe62069f0ba9019f0725f54b;
mem[704] = 144'hff0ef463f96ef7d60374f34a0b9e06080d65;
mem[705] = 144'hf5ec06e8f4df0ac5f5c00d130bdcf7e7fb58;
mem[706] = 144'h08540183f51af1e6042400d10be80aedffb3;
mem[707] = 144'hf3c900f7f6e70e76eff603e1f941031a00eb;
mem[708] = 144'h01d4f04109440061f07e020d052bf36af76d;
mem[709] = 144'hfcb1f00bffcbfff104a5fb80fa94f0b306c8;
mem[710] = 144'hf50ffd6b03f1f8e5f1740907ff9002db0852;
mem[711] = 144'hf8cbfc40f3a000be0cd5f687fffa059df1ab;
mem[712] = 144'hf4bd0e86ff7b0b2f03ad01f200b1f6b7fd26;
mem[713] = 144'hfbd00596fbe5f2f5f6c4fca1f9130cda0bb2;
mem[714] = 144'h0ddaf8a808b9f7e70736fc1bfffcf14f013b;
mem[715] = 144'h0563febbf5b7012a0becf012f635f150fb75;
mem[716] = 144'hfab505860b7104d505b20f78f81b0945f354;
mem[717] = 144'hfb5df911008409fc0902f2dafe4a08ad050f;
mem[718] = 144'hf645fb87f566ff1c0f850b50f237fee4fbdb;
mem[719] = 144'hf39a04140cc2f7a10359f805f0120a68f7f3;
mem[720] = 144'hf89cfc43f262fc1cf074f78efc2e0b4df2df;
mem[721] = 144'h0899ffa20c59f705f40b0aaa0f1df942025a;
mem[722] = 144'hfeb3fdbc08f3febb0d920a820b0ffc350326;
mem[723] = 144'h0f1bff5e002806b8f6c6fee6f640f7bcf7b1;
mem[724] = 144'hf2f2fcbc078af1ca06a9fce30481ff96f479;
mem[725] = 144'h019ef0da0d70ffe9f3b70d5ffa430f88f0ff;
mem[726] = 144'hfbc608400959f235f05cf05ff5b00c9e0529;
mem[727] = 144'h0e08fd90fbfaff21f031f5f2fa59072602c8;
mem[728] = 144'hefa70c92f4bfff8bfd04035ef866f90c00de;
mem[729] = 144'hfd04f7a90ab7fc7ff7b20836f0c0f4aef191;
mem[730] = 144'h07faf39ef9d1f669f5e1f53a08980e4a0680;
mem[731] = 144'hfac0f2e4fdc1fc35f4570fedf86df04ef3ac;
mem[732] = 144'hfacdf433faf00a330ed5f8eb04bf0781004f;
mem[733] = 144'hf465ffdef2b10baaf670f876f499026ef10e;
mem[734] = 144'h0f28014cf4d8f3ecfbc801fcfee9f2fbfaa0;
mem[735] = 144'hf9c606c906690fc102a90de2f999f4a80cd8;
mem[736] = 144'h086a01fff964f896faf00f1707f7fef7f831;
mem[737] = 144'h0cb9f276f0e60995f053fc5bf3bef09cfe9d;
mem[738] = 144'hfc49fcbcf5a4fa300fdcf36b04bcfe7ffba9;
mem[739] = 144'hf3e0f974f7d10cc4051109fdf4feefccfb6c;
mem[740] = 144'h0740f9f80ed10a9ef762f2bb0b2cfee1037c;
mem[741] = 144'h090d0e1ff7740636065f060e021201e7080c;
mem[742] = 144'h0772fa53012305130a180592f5a107c50381;
mem[743] = 144'hf53ef21efda0088a02c2f97b047f0b3f035f;
mem[744] = 144'h04f5fa4408fe0504fb4100a00045f652fbbf;
mem[745] = 144'hf61ff3690c8ff1c90e340e0200acf9dc0df4;
mem[746] = 144'hfabeff6df5e7f8db0c4c00140b780752fbab;
mem[747] = 144'h0aeaf408f29bf802f0460e0d0ecdf04a0057;
mem[748] = 144'hf93306f106f202b803180b8dfce90174fc3a;
mem[749] = 144'h091ff60bfc4b0e89f0e5f4a905c904070cca;
mem[750] = 144'h03e5fcf3f087f25f0f07f3b70d3c0f660563;
mem[751] = 144'hf5d1fb72fe44093702170bb90e98f01bfdeb;
mem[752] = 144'h08b50448f782f6e60113065df503feabfdaa;
mem[753] = 144'h009500f6f3b6f7f40818077c0044fb1d0aad;
mem[754] = 144'hf370f20609c40d20f4cd03bf0728f25d0608;
mem[755] = 144'h0cdaf482f084074af438fb9af97908840b30;
mem[756] = 144'hfd71fb00f38e080afd0001600bf401220b7a;
mem[757] = 144'hf885fbf20d78012af34b0fb306050a16f5db;
mem[758] = 144'hf0f5f04ef7f904180ab50cbf0320070bf610;
mem[759] = 144'h099af1e0f65c05a9f50efb3d086d0b17fadd;
mem[760] = 144'hf4ae0170f809fdc2f06a04900ba40af7f3c8;
mem[761] = 144'h0164f33802ed0896f171069d00a9fe07fbbc;
mem[762] = 144'h091209bb0da10e8b05c6f4a6f34efeb8f316;
mem[763] = 144'h071bf6d1088105bf064802a5f825f332031e;
mem[764] = 144'h063701b2f04f01a5f64ffbd3f89700c30505;
mem[765] = 144'hf4c10a33f0a1072ffb420fa40e8f0ad609da;
mem[766] = 144'hf38df25e0238ff26f46a0137003e01c4f296;
mem[767] = 144'hf2f10422ff7a0b0aff54f707fe7b0a5afbc3;
mem[768] = 144'hf0ae00b1fa7f043a0414051af1cb0981027c;
mem[769] = 144'h0b04053df7fb0fe50004f947082cf4830a11;
mem[770] = 144'hfe54069e01fb0cbbf0ca0223f879f0ce0b6b;
mem[771] = 144'hf278fa680e2eff11059104eaf796fcac0a9c;
mem[772] = 144'h0525f5f8052ef4ba08f2fd1a0dee0cc50b91;
mem[773] = 144'hfb08017cf4460cbd017a0e95034bf9be028b;
mem[774] = 144'h01e20c1e0c6ff2cef5690eb50e95f3e4fd40;
mem[775] = 144'hfcaa0a9ef920053dfab6095cfcadf7bbf620;
mem[776] = 144'hf53a08d1f455f6da0e19f8ad0df1f26e0eb1;
mem[777] = 144'hfa8f02110352f6df09ed0788087bf0810fb9;
mem[778] = 144'hf62a0dee01effbc3f3c2fb32009b015f043c;
mem[779] = 144'h0f03f7c5fdfa06db011dfbfaf1c9041f027e;
mem[780] = 144'h07b0ffb8fe23fb7a0c5dfbb6ffa8fac10455;
mem[781] = 144'hf8d80f9afab1067f0e9903a909bb01b40c8e;
mem[782] = 144'h01360702097ff08208480acf0eadffa6fd71;
mem[783] = 144'hf14204d9fad3090cf830f172fcea011a08fc;
mem[784] = 144'h0c21f9c40afb0994fe4bfa6dfad90a470cc6;
mem[785] = 144'hf74d035c08420df906fdf940f384fd1cfa50;
mem[786] = 144'hf49c06efff0a04d60d29f859f3e20ec10cd2;
mem[787] = 144'h0b9d0a180bc80397fba8fac2f69a0f05f1af;
mem[788] = 144'h099afc45045c098d012003ae09bdf13ef445;
mem[789] = 144'hf34f01aef6d20deb06f1f27b0d21f2fe029f;
mem[790] = 144'hf6b00c590afe050f08f4f7570d6d087e0e45;
mem[791] = 144'h000bf3460db6fa96fbb1f1390169fe2cfac3;
mem[792] = 144'hf8290607f965f981f467fa010b1ef5670818;
mem[793] = 144'hf12d066a032a0cea093807fd046af645013a;
mem[794] = 144'h089bfc4ff692f71f0527f00c0fbd07120044;
mem[795] = 144'h01a4f794f3d9f89ef64bfc7ffa59f155f786;
mem[796] = 144'hf30108450d36f1ca030cf671f81afb3f02e7;
mem[797] = 144'hf8da09f804ecfd08f707fe2e0e7e0aaff072;
mem[798] = 144'hfc93fc7ef18a0503082a0191faaff46b0ad9;
mem[799] = 144'hfdb2f2bf02ebf95afd7a0ce205290d300168;
mem[800] = 144'h0956f1c4f19af5a409a9f0950a0ef3edf635;
mem[801] = 144'hfdaffc980bcf008d0790f97bf106f43dfda2;
mem[802] = 144'hf87e043cfaddf7d6f4b7f011f466f4450e5f;
mem[803] = 144'h032a02a90c63fd1df99ff3b70067f0060c4f;
mem[804] = 144'h0854e7a1ee02e742fbc6f27cf090ecb5fdfb;
mem[805] = 144'hfdf8f80a0855024f09fef92bf8eeef59097e;
mem[806] = 144'h0d41f23101d2f319f932fc1101860252f393;
mem[807] = 144'hefc2ec4ff2bb008c0116ed41f092f50bed83;
mem[808] = 144'heb79f5d2fcbf0411f2910466e9fef713f5c2;
mem[809] = 144'hed51ffb30cd9f6e2f7a2f0a00c3f0da5097d;
mem[810] = 144'h0632ee7cf4950908091bf7ed05e5eef6f56a;
mem[811] = 144'hfd09ff3cf82df062f0c601f506e40ce303d0;
mem[812] = 144'h0871f73007aef127f3cdf7c70850fc4cf993;
mem[813] = 144'h07cb02370cf90855f473f3240038004f0aa8;
mem[814] = 144'h06a40400f8a00809fe74fe37fde8ff55f28d;
mem[815] = 144'hfd01f390f4d00ecc001d0ae1f72ff02bfc26;
mem[816] = 144'hfa51f47af4ce0c95f4950234fc08f0a60eba;
mem[817] = 144'hfbbaf356f6bf0cb4f858f097fe140a3b053f;
mem[818] = 144'hfbf905dbfbdcf772f2def93105530dc40ccb;
mem[819] = 144'h0a4ff6ba0935fb840d4efdcaf967f2ceeef4;
mem[820] = 144'h050b0d1ef981eee1f79a0239f95107a307ff;
mem[821] = 144'h087fffed07dd05b20aaa001ffc770ae509f0;
mem[822] = 144'h00140761f12f03870d48022ef8b90f2a0197;
mem[823] = 144'hf01f014d03d6fe67f9f9f35b01e604dcf3a5;
mem[824] = 144'h01810c8df23008cff8f60822f64af4bf0acb;
mem[825] = 144'hf5fdf18b0a2d007dfaf309b203e6f2ab089d;
mem[826] = 144'hf9df0849f9f9fc900251feaa067cefcf0831;
mem[827] = 144'hfc19f0c5020d056a0c5e0f24f145fc2ff012;
mem[828] = 144'hf7aa024f080406dbfa170a33f3dc095dfb6d;
mem[829] = 144'hf3470bbdf47fefa404cbfde9f8c800eb0b35;
mem[830] = 144'hfa8aff5dfb37f43cf9430d8df7f20c40f6b1;
mem[831] = 144'hef40f44d0def0ef1079801dcf989fa88fe2e;
mem[832] = 144'h0555f419ffdf07a50f25f1240f09f194fdb5;
mem[833] = 144'h063709ea053a03ebf5ee0d4df415078802e4;
mem[834] = 144'h0d66f80ffc21018b06e60a47faa8f775f01f;
mem[835] = 144'h06d2fefafb80f7e9f226f0f3f8dc0e74f1d9;
mem[836] = 144'h0a3cf077fb9e060ff8200e3bf314ff5808f7;
mem[837] = 144'h0c5efb4c05affd23fb40f1edfa43f1ecf439;
mem[838] = 144'hf4e8f065ff99f5430be60a00f6e6f022f13f;
mem[839] = 144'hf540efeef506fa87f723ee86f32806c5f099;
mem[840] = 144'hf3c004c4036ef99d0c2903b10ea2f077f3b7;
mem[841] = 144'h05c3f6a60a0bfad1fd6604e00011001a0497;
mem[842] = 144'h00e7f3580bfcf91c01ec044105590751fa2a;
mem[843] = 144'hf64207030e89fd7e0df40437011df92f0c2e;
mem[844] = 144'h0018f45c021c08530325f01afd89095cf838;
mem[845] = 144'h0f1d06b0fa330070efad04c106aa0d20fb99;
mem[846] = 144'hf4a1fb1b0581f45003820f9b0f4707cf0b99;
mem[847] = 144'h0949f604f5d8f607f869fc7ff009f6370782;
mem[848] = 144'hf979068402db01190a89f86b035cf43e08f5;
mem[849] = 144'h0e35f7d109eb087ef1d805ba0f14f2fbf3ee;
mem[850] = 144'hf5fdef87f81efc75f5980ca4037ef231f150;
mem[851] = 144'h0e960f34f1f00af3f7700101f1ff0b31071b;
mem[852] = 144'h0eb4001e01b20bbaf78705b90631fb9a07b0;
mem[853] = 144'hf3a80a060a25ef62059d05a4f6b2ff2f06cc;
mem[854] = 144'h0a51f24a07b1f947f62f0bdc081709c5f5cc;
mem[855] = 144'h021a0753085c0641075500a2006100fe0467;
mem[856] = 144'hf91dfe90f41c0d89f2defdc7fd72f4bcfa30;
mem[857] = 144'h09890337fe1fff6609490e380294009af24a;
mem[858] = 144'hfede02ef0685fd02f7e8fd9802cef9f0f2d7;
mem[859] = 144'hfddb0b480528faaf0f2608eb0272ff0a011e;
mem[860] = 144'hf834011e0e83f582f22205f202be02f0f1e9;
mem[861] = 144'hfea004d6f0010a9807680d010d2ef166fe7e;
mem[862] = 144'h0b30ffcf0c6508a3f9a3fe6c023208e40a24;
mem[863] = 144'hf7780aa1f01f058bf21efeae0cca03bff056;
mem[864] = 144'h0d05fbabf3d00dcefa76f604faa3f5000077;
mem[865] = 144'hf6a8ff980d67014dfcf5f7500dfa0924ef5e;
mem[866] = 144'h0426fad00f0d081df51b0fdc08c405710bc3;
mem[867] = 144'hf50005dd05640b07fbcb0dac0aa3f63af9f6;
mem[868] = 144'h04aef518efd3fc6fffdf031efdc8f1320975;
mem[869] = 144'hf459ff2cf1edfef9f9d7f913fbadf4850a2a;
mem[870] = 144'h073af8380b97f9d50107f4fff592f3c6ffce;
mem[871] = 144'hfa43fb4701b502e6ef5e0544087e00daff4a;
mem[872] = 144'hf4a1e876e5a1ff1cead2e7e5f6e5f932fbfa;
mem[873] = 144'h066e0a6cf385f89a01b9093c0c88fe42f2a0;
mem[874] = 144'hfd22ffb7005d041d0bdd0d14fd86f4490c2e;
mem[875] = 144'hf8baf57cffcdf26af2e10dfaf2f1fd64fce8;
mem[876] = 144'hf38500820aaff0310a0af46107450ea8f153;
mem[877] = 144'hfa93f44008dd026cf4d3f173fea0f3a105f1;
mem[878] = 144'h028dfbdefb59f16c03b8fd650ee20d210231;
mem[879] = 144'heffc0000fde9fcc7038202ccfa660209fef6;
mem[880] = 144'hf8ecf37d043d01ca0376fe570db003f0fa80;
mem[881] = 144'h0809097c0b9cf5f30626ffa60dd0f6daf3b4;
mem[882] = 144'hfc770cad0522fc58ff52f045076ef2acfe2f;
mem[883] = 144'hf143efd60478fdac0533f4d4f36aff97f563;
mem[884] = 144'h023cf17ef3b60913f6410c22fae60389fad9;
mem[885] = 144'hf8fbf329f433f580fd55f2ce0dabf2170d1e;
mem[886] = 144'hfa5a04f4f2120aad06d10113fda90da2fcf7;
mem[887] = 144'h0c7af671058c00490dd5f8210baaf547ee8d;
mem[888] = 144'hef4c0b6f07c80971f085f3d301e2062bf717;
mem[889] = 144'h090706000543f3f5f4b70b56f2ee0c71fd85;
mem[890] = 144'hf2c9f75ff1cbf4e907a80731f48cf75d063b;
mem[891] = 144'h085d0e8506fcf6b30193f4150e01f17005e0;
mem[892] = 144'h0314f3c4effd035bf308fac6fdc0f5060471;
mem[893] = 144'hf219fbb1f9bd03ba078206a3036ff76ef455;
mem[894] = 144'h09be03360e98fc37f3dd02f9fd5af707f199;
mem[895] = 144'h0c42fd5ef973f77afde204f2fcd80bc1fc92;
mem[896] = 144'hf55a06360af4f6e5f9b208940cbef0ecfdc7;
mem[897] = 144'h009f0035fc820ccc0f25093f0f79f35ff6ff;
mem[898] = 144'hf60907c0002af87e0e5b0773078ef1fdfe29;
mem[899] = 144'hf24b008afc5efbc10681f0a704dcf1b0095c;
mem[900] = 144'h0e3cf6780b3af9a0fffd0cef09bcf7bf09ce;
mem[901] = 144'hff100625f5dcf564f68d0d31f551f1a1fb24;
mem[902] = 144'h03baf991ffcff6ce096cf0f0faf2fa870cff;
mem[903] = 144'hf1fff23c05f1f0a4f8caee440667f45902f4;
mem[904] = 144'h0014fa380083f2d10980076c0bb8fd440b87;
mem[905] = 144'h0cf6fc73f29ff92b0a560d1ff85cfa520893;
mem[906] = 144'hf90cf9c7f1b10bd6f7f50d6efb4b02e8fb75;
mem[907] = 144'hfc95fa5f027df31ffdf704ed06820c55fe66;
mem[908] = 144'hfdf7027ef84901beff7009b5fed1016504e9;
mem[909] = 144'hf0040070006ffade059006c9010d0c85fc93;
mem[910] = 144'hfbdef47d0feaf7980fc5fad7f5e502dffc3f;
mem[911] = 144'h07dafd550c34fda6000efc6afc1bfceaf759;
mem[912] = 144'h07ccf56908eb0b3bf2cf04180b33feff06f7;
mem[913] = 144'h0849f9800dd1001b0182fc2406260505fe18;
mem[914] = 144'hf0f4f954f655fb1907b6f2b5f1df063efa93;
mem[915] = 144'h0e5c03d0f3740038f070fdf1efb403c80aa1;
mem[916] = 144'hf6b1fb85fa37f865f8ffff83f1b7003a0361;
mem[917] = 144'hf6b0f27f00b60e1f0265f62c0340f7c3f229;
mem[918] = 144'h0370f139f06409d20b100300fd42032a033f;
mem[919] = 144'hf82cf217f1a6f3a2f357fb64057e03690c67;
mem[920] = 144'hfb9bfa390634f67309affdb2fc42fa40fd7b;
mem[921] = 144'hf6ddf4c0f1d4f21e0bcbfa5bfa6a0ce9f833;
mem[922] = 144'hf48a0cb4fdff06d0f4c903f4f68e097efefc;
mem[923] = 144'h0fcff0aef04900af012807f8fe360f9dfe3b;
mem[924] = 144'h00c406f0f1130e0ef5f80a77fdc106ea0c8a;
mem[925] = 144'hfffd0537fef5f79bf72b02340692fe8b0757;
mem[926] = 144'h049c0326ffa40eadfbc2fe02f8840cbbf166;
mem[927] = 144'hfde7f3c20700079708a0023aefaff914f4f8;
mem[928] = 144'hff0b0958f85d0b8c00a4fa07f82605a20d44;
mem[929] = 144'h0c0d0b73fdea0faef11cf6e3066f0e6b00fe;
mem[930] = 144'h0988f5b0f3340de505830444f73ceff30df2;
mem[931] = 144'h0ea1fb57f8a707fa0805fc690c0b02be07a0;
mem[932] = 144'hf63efcebf15a0395f78ef561f5cff06df577;
mem[933] = 144'hfb14f7b90b3f06ffef41ef4bf420021ff56b;
mem[934] = 144'h03480525f5bb01bbfeaa0c4d0973f1b4fb7a;
mem[935] = 144'hfeccef7cf83bf8de06b303eafdd00a6403b4;
mem[936] = 144'h00c0f626f352ff0afadb0617fdeafef707c5;
mem[937] = 144'hf11ef41b05a60199f2c7f9590573fc77fa1f;
mem[938] = 144'hffe700410163f5060131f2fcf65c0350f615;
mem[939] = 144'hff6100f0fc26ef8d081408ca04cbf42c0b78;
mem[940] = 144'hfd3e0d70032c08eef2910ed4fe6df127f617;
mem[941] = 144'hfe27081908460b0f0257f1520575ff69fe60;
mem[942] = 144'hffd90914008cfc960306f2440e3ff9a6fcba;
mem[943] = 144'h04c6f4030f49f21c0c7a03c902590041fe39;
mem[944] = 144'h04e80070fa10fa040a67f958f922f39d0c73;
mem[945] = 144'hf799f1c1f513fc0202980703fbe109ef0f8e;
mem[946] = 144'hf9fbf5360c6dfbedf23f09c3fee7f50406ce;
mem[947] = 144'h0dc2f7fe0592f1c6f9ff0edaffcd059ffafb;
mem[948] = 144'h0f640879f603f174f7fe09f3f8d60e81fba0;
mem[949] = 144'hfc0cf3050290f7a7fcda0ba1f806f8bdfb66;
mem[950] = 144'h02e70231fbd002b00b80ff40f0cf094ff1c4;
mem[951] = 144'h04a3081efdf70b3e0df0f381f254f70deff1;
mem[952] = 144'h046bf1d6fbfb0d2c0fb60e7feff9efbe0bd3;
mem[953] = 144'hf667048d00810142f3170bc408ea07bf0d0d;
mem[954] = 144'h037209d8f0daf2a70a7307c90649fc690bab;
mem[955] = 144'hfef7fa680052f6adfcaef29cfc3506590f2d;
mem[956] = 144'h09a709eb04e10410fc2804c4fd670c88fb28;
mem[957] = 144'h0e21f8ddfe59f6e2f83607e1f448f1240532;
mem[958] = 144'h0fad074d063e08e60ed1f5b6f21bfbe7f8b1;
mem[959] = 144'hf9ac08b205220cabf8b7fdb4f4dfff480795;
mem[960] = 144'h0ee7011ef5c8fa6b0858f27608e1f72cf420;
mem[961] = 144'h0e0d072df9cdf66ef89f08a4f20903c906b5;
mem[962] = 144'h07e2f26cfb9aff70f9cb0a8f0cc0f8c60e08;
mem[963] = 144'h055200f4ff4bfe8cfcb5050e0d410a690e6c;
mem[964] = 144'hffe30a64ff3ffa61ff50f0b907b40cde05f8;
mem[965] = 144'h071cfbfff9d3f2c2fbfe055a0926f70d0d1f;
mem[966] = 144'hf05ff50b069b04ac03fef83af6b6f884011b;
mem[967] = 144'hff4bf1a500690879fbcef6e50bfe0a14f09b;
mem[968] = 144'hf1900cfc021302a0f85df7b70f02f0ebf677;
mem[969] = 144'h0ec5f0bf0ce7f05f05b7ff9df7140f2cfeec;
mem[970] = 144'hfd2602680570f3b5f730f2dbf53602330c65;
mem[971] = 144'hf6d3f7b5f0ecfaabf99efa56f51505aa02ef;
mem[972] = 144'h04affd2000e90f400e37f900f84df9faf4fa;
mem[973] = 144'hf18b0f0703ba05fafe47009506570beb0080;
mem[974] = 144'h06ecfb750552fe07f1ca0f070f5b0289ffaf;
mem[975] = 144'h02d00ec304f5fb30f1bbf59d0e97f7a00d5c;
mem[976] = 144'hf984f5c2fdf80ad10e49f57d065df911f3cc;
mem[977] = 144'hf0bd0c99059006fa012205f3fe20fa5e0f1f;
mem[978] = 144'h0267fd94fe75f79d0dfa0226015af9fb00f2;
mem[979] = 144'hf3f1076606b507b5f24706a0ef550741f91b;
mem[980] = 144'hf68a0d07fba50af7013bf32efca4ffb6efc0;
mem[981] = 144'h094e048705ac0fa6f3f4f4cef6fdf62dfd9a;
mem[982] = 144'hfc0800c6044bf4f7f6c6f58d0bf5f0360066;
mem[983] = 144'hf203fe51fd0504b704f6f5600a23f2eafc5b;
mem[984] = 144'h08a5f8890330f7b0ff31f31c0c72fb40097f;
mem[985] = 144'h0ccafc5efe570b5ef1890954f785fd5ff659;
mem[986] = 144'h095ef9d907330f7df2a5fdcbfeb1f1280ed6;
mem[987] = 144'h01b8f21aff50f0ed013f014401210cfd034f;
mem[988] = 144'h0f5bfc14eff9fdbf008ef098fb10012b0b71;
mem[989] = 144'hf10b0ef609b1fe630364f1630280fc8ff349;
mem[990] = 144'h04850c2503100eba022001b30eb00dfa0f1c;
mem[991] = 144'h04abfd76f54100ec0d4208d604250e2c0d0c;
mem[992] = 144'hf23d086bf9c8ffa0fa860701ff84f4dc0bfa;
mem[993] = 144'h01d2fe950d91f932fdb703ae0151f892f163;
mem[994] = 144'hf942f854f13b00f00b6bf852f1bd063defd1;
mem[995] = 144'h046df22303df05d1f9b9f24b0566f0ce00f8;
mem[996] = 144'hfb65f10609d8fc58efe90be1f96000e7f48a;
mem[997] = 144'h072e0c2feff903590663f4ddfaf4f86ff8c4;
mem[998] = 144'h0df00dd30ee2fd48f3d20b9d09fd097f0c63;
mem[999] = 144'h0b8b07b1f41af9ccf73cf547f2e700e7f212;
mem[1000] = 144'hf05d0a2ff4cffbf30846fb8ffcee048c088c;
mem[1001] = 144'h02a3044d05ecfc9dfba609640d5f01990a55;
mem[1002] = 144'hf669f0850d780364f7060f5009bffef707fb;
mem[1003] = 144'hff37f2860da60de0fce002330be7f8d605e4;
mem[1004] = 144'hfcf8f9f4f7290e0604c4012001b20cc1f8d2;
mem[1005] = 144'hf8a90b0ffc28f5cc016205370495f6c40bcc;
mem[1006] = 144'h0a670449fc73fe850eb2fec8f047efe302cb;
mem[1007] = 144'h0e0fff2305500a190ab60091003cf586f01f;
mem[1008] = 144'h095200ccf8f0f1a8fc78f2dc0ef7fa5504e2;
mem[1009] = 144'h0c7efed70de7f33ef396085e0149fde5043c;
mem[1010] = 144'h0a17f7950b39f6b90c81091a096902480a3d;
mem[1011] = 144'hfcabfbe9f0a403b3f311ff0b08bdf1cff5f1;
mem[1012] = 144'hf6bdf57cf62ffe91ef8cf7e0fdfd0aa50276;
mem[1013] = 144'hf59ef758f8b2fe62f9a80bb5f94e0d22fdde;
mem[1014] = 144'h04d40dadfbfffb1ff4760d430a86086106ef;
mem[1015] = 144'hf9520067f99d0c90f55dff9af7430986f6fe;
mem[1016] = 144'hf1f4f61d07f5f51ef515f744eea8028ef482;
mem[1017] = 144'h0d0a0dc0fbeff717f89900eb0c26f24a0305;
mem[1018] = 144'hf633f4610462f88d0fa80c8f0b55f01c098f;
mem[1019] = 144'h05ba002df6e205c600d20c18fc4efe4aefb2;
mem[1020] = 144'hf90f017ff5fefe6e0ca404c30502fb3afd00;
mem[1021] = 144'h002d0b42073f0a2ef90bf16500a3fe600de7;
mem[1022] = 144'hfc0dfdfefc42f8cf06f8fc5a0e740c2ff263;
mem[1023] = 144'h0b750e71f698016f026b0e9efaaf00190b58;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule