`timescale 1ns/1ns

module wt_mem7 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h06d70204f94b0d0ff51a0c270ed7f501f8cc;
mem[1] = 144'hf50f026e04b10c82f587fc1403000c23016a;
mem[2] = 144'h0172f682f72703c2f9720ada02a0feebf60e;
mem[3] = 144'hf63affe10375f0dcff3a03b007ad0cc90b48;
mem[4] = 144'h063a0615f3e3050205220fce00eef58af549;
mem[5] = 144'hf84bfddf0bd5f4b400b00062f8c7fe730e02;
mem[6] = 144'hfceaf7d7010f0a9e03590b990a6b025df83b;
mem[7] = 144'h07ed0929056ffbd70e28fdebf6b3fa400a71;
mem[8] = 144'hf68ff0ddf15a01800386ff7703f5fb74f602;
mem[9] = 144'h012cf90f08420673fd140a020fd8fec2f2fd;
mem[10] = 144'hf1f70373f41608f607b70194faccf359ff86;
mem[11] = 144'hff8cf8a4fda10899f124fe73fca9058b0383;
mem[12] = 144'h078bf3c7f9f7fd5cf08e04c1fd84f9110e87;
mem[13] = 144'h0bb40fd503230417f716fc35fb4104cff45e;
mem[14] = 144'h0577fa9bf95b0f61051c05b70844f7af00c4;
mem[15] = 144'h09eaf45f0d4dff63fc7106b70c660d720395;
mem[16] = 144'hf09904f4f3ebf2bcf75ff85f0f4ffcbef7fd;
mem[17] = 144'h00860a5402bdfbd70af20bb50dc9fbb40dd2;
mem[18] = 144'hfc7b0e020a55002906aff42404b5fc7df1e0;
mem[19] = 144'hfc44f16cf08002b6f7420ba3fe940aa7f25f;
mem[20] = 144'hfdb0fd720689f811f3a3f7c5f94dffa50916;
mem[21] = 144'h0dc2f58ef00509f7fb52fa0c0713f5d90645;
mem[22] = 144'h0251049b0f0af1fbf7070b02ffcc0ab2000d;
mem[23] = 144'hff36f0fffe5e0cedf18cfc09019409a20913;
mem[24] = 144'hf072ff1b04f20988f7e5f528f463fb77f8c6;
mem[25] = 144'hf4f5fd9bf59106ae0c1004360240fc7103f2;
mem[26] = 144'hfc99f506fa02fc0ff5e40874035ef30bf754;
mem[27] = 144'h0d78f502ffd9f1980ac90fc402e2f53afb24;
mem[28] = 144'hf47afdf9f96f03960abaff29f81ff5fcfa7a;
mem[29] = 144'h03ee0312f0e7f72f02f900350252fe1cfccf;
mem[30] = 144'hf9b60940fa42f513f8d30a910b62f77c0a56;
mem[31] = 144'hf45bf7870b49093df7bc0620f2f8f3480743;
mem[32] = 144'hf50201ad0d1bf0170c05f46af91df1790ad1;
mem[33] = 144'h0be0f0fbf6e0f2a9081a05c1fec3066201d1;
mem[34] = 144'h09dff29afd8defd0f82cfaeaefe1f090014c;
mem[35] = 144'hf2d602b0fddefb1a0558f47102c704a107fd;
mem[36] = 144'hf57df87e06acf5fc01a1058003790dca0e72;
mem[37] = 144'hfd09f40bf87dffd80b9e0ba2f3c70313f1bf;
mem[38] = 144'hffc70d97f777ff51fc2505b0ffcaf39e0ab1;
mem[39] = 144'hf3dbfd2b0512f553ff81f053eff8f4fef3ab;
mem[40] = 144'hf18afbf90c4900ae09b6069ff389f77dfbf7;
mem[41] = 144'h0c76ffa9f909feb2f1f7f86701bd0c8c02fa;
mem[42] = 144'hfc9bff8cf5b7ff3ef88a0b5d01f20f9af0d2;
mem[43] = 144'h09c5f1800022f5e00345f0abf7bd08bb0f81;
mem[44] = 144'h03f20209052cfb050b830cc0fab0f669f661;
mem[45] = 144'h06f601e40e01039709f00bca090c02710025;
mem[46] = 144'h062c0c93f902efecf9e1f367fbbe02d8fbe5;
mem[47] = 144'h0a45f163f9ed0dab01ffff79fca107a7f6cd;
mem[48] = 144'hf8410a4a0677f64809aa0b300321093108a4;
mem[49] = 144'hfb7cfaf3f69106f40e8708790b310e40038f;
mem[50] = 144'hf2a30ce2f98e00650709061a0ab3fc270c1f;
mem[51] = 144'h03c700e2fb7af0bcfa4df433fa1403180d1e;
mem[52] = 144'h0e9606d6f260fe0a0585f882032ff6a00b7a;
mem[53] = 144'h026700c0f485ff1ff71104d409b206a30441;
mem[54] = 144'h0d61f40a0a99ffa0082df8440a9f0d8cf6c4;
mem[55] = 144'h0d4ef820081ffa130bf5f0d50b3ef5d6045a;
mem[56] = 144'hf5ebf5c60ac605d8f15ef38df1790c3dfcea;
mem[57] = 144'h045304cefaa6fc39fc030d2b0866f95dfe60;
mem[58] = 144'hfaa2fea2055408def3f40a6fff570c1d04b2;
mem[59] = 144'hf339fbf9f8d8ff3e0c23f14bfd2bfd36f6c4;
mem[60] = 144'hf29cf3b3f0620e36f0520468f057f6c60073;
mem[61] = 144'h0d91059efcb900b80d5ff9e303e7f4c40629;
mem[62] = 144'hf4b2f1bc0757f602fc4cf3290943f98c0950;
mem[63] = 144'h0ac7f2c908e6f95f098403e9f0dc06be0a69;
mem[64] = 144'h01cb0be30b0d05b10e160d15f2e2f2f0f058;
mem[65] = 144'hfd01f453fffcfb8b0cdc091408ecf94005ae;
mem[66] = 144'hf7affd8af5c6f03d09abfbe409c307bbff1b;
mem[67] = 144'hf69af63ef1a1fb8fff6b01cbf6050909f546;
mem[68] = 144'h06bb035efa7cf4dd0040f7120bd40d760251;
mem[69] = 144'hf63befe5fbacf5f9f7ee03d500e0017a0ec4;
mem[70] = 144'hfdfa012107a9ff92f5ea00890eb00a64099e;
mem[71] = 144'hff20f43fffb6f7310a6e0f5cfbe4fefe07d2;
mem[72] = 144'hfad10069007803290502f68506930028068d;
mem[73] = 144'hfc7b0716fef5f13f04e1f0560e0604bff119;
mem[74] = 144'hfd79fa870f55fa8a095cf741fd92051a09e1;
mem[75] = 144'hfb990a30f0670509f7ef0e1003f20be006ac;
mem[76] = 144'hf2910909f0cf0c06035f09b00cfafe8bf3d5;
mem[77] = 144'h0906013506620a510afff767fac2f8d6ffce;
mem[78] = 144'hf7730ad80d060e7b015d0cd50c92fc1a0f0a;
mem[79] = 144'h02ae06230d3ef667088f0f51f421f2c8fb30;
mem[80] = 144'h0a830a580238f919f92e0619f395fdfbf0c0;
mem[81] = 144'h0087015a02350e1df4fd02c1f0b80ac0f7fa;
mem[82] = 144'hf0d303a9f6aefbed0016f4df0c2df49ef366;
mem[83] = 144'hf30ff98ffa16f52ef4ea07c6f671f00e0015;
mem[84] = 144'h0f6308bdf0c20915fa6dfc3cf5020fbc0fb3;
mem[85] = 144'h0dfa07310819f35a02fe09c0f314f7670373;
mem[86] = 144'hf7c1046cf0b20f640881f871fd450275ffdc;
mem[87] = 144'hff3fff6009a3f160fa0ff5b90a68f82901f4;
mem[88] = 144'h018806590ca7f1a50ce80ee2f7bef9c008ec;
mem[89] = 144'hf7edfc87f414f713f90704e5f06e0cd5f2d0;
mem[90] = 144'hf996f6f3f9f2003f03c00272f7880ba2f131;
mem[91] = 144'h022b07c60cb40444f5e70960f0e802e8f708;
mem[92] = 144'hf2ab09dafe25f3fcff3bf75ef21e0eacf74d;
mem[93] = 144'hf549071fff22058cf9810ddafe71092c000a;
mem[94] = 144'hffde0083f09afabe095f09210bbdf6a5f727;
mem[95] = 144'hf1e701730910fdeb00b8fdd401a501f201a6;
mem[96] = 144'hf97ff368f04ef90efa3b0191fea7fb0b00e2;
mem[97] = 144'h0a8309c70303f3da0b4d060bf865096400a4;
mem[98] = 144'h0b14fe1700f80939fdb8fb39f4f8f20e0c41;
mem[99] = 144'hf1cf0f37fa0c0c97f9de004a030afc4200fa;
mem[100] = 144'h0ec5fc57f03a0099fe8b0cc80cf801c0f1be;
mem[101] = 144'hf86903ca03930e17f55df0f70d1aeff70522;
mem[102] = 144'h09bcf11a04910e1d038b039f0d1dff870b8f;
mem[103] = 144'hfbfbf1fdfdbaf9730153fde4ff5e01b1f4a5;
mem[104] = 144'hf28108a6f70b0647f67a009dffab030efa62;
mem[105] = 144'hf43c023af065f941fcabfcc0fe2d0f550941;
mem[106] = 144'h086ff011f759f10101fffcf503fbff8b0f02;
mem[107] = 144'hf88cffaa074902b6ff07fac8ff1ff6c2fd6f;
mem[108] = 144'hfba9f5d7062307a8063c0e14fb560cc909d6;
mem[109] = 144'h09480403f2dd038c0d20f8d9fa000848035f;
mem[110] = 144'hf796f91b07ec000606320fd5030202910df3;
mem[111] = 144'h0a42f7a7009df52b08edf8d5f02eff670c38;
mem[112] = 144'h0933f714f46e0baef0990188f606080100c8;
mem[113] = 144'hfd6c0b23f9ac06d8f09400dbfac700b50120;
mem[114] = 144'hf041f04ff2b2fe3006ad048bf2af00e0fe12;
mem[115] = 144'hf0d2f517ff9cfdf1f413f3c9f75f057903f7;
mem[116] = 144'hfcddf68609b6fd32f96ef3f1f77b0244f2b8;
mem[117] = 144'hf138fbbff76df41605320c1d070801340d72;
mem[118] = 144'hfe080ded0c4df4c606fbfd280112f75fffdd;
mem[119] = 144'h0fd90bc20360fef4f1eafd290bb50eae0411;
mem[120] = 144'hfaff052cfe2808b1f40504de019500020e30;
mem[121] = 144'h0a58fc29fd0ff1070337fd6001a20117f1c7;
mem[122] = 144'h0a8cf02fff8b08dd0aa8f519f254fd780a40;
mem[123] = 144'hf8dc023af8b5f143f5d6f019ffb9ff51f8e4;
mem[124] = 144'h0e2df55ffa2af8cefd80f555f8750d71fb36;
mem[125] = 144'h0009f6c6fb8e0552f96506c7f308f2bc089e;
mem[126] = 144'h06ca0b66f284f1ea01520daa08dff86cf2c6;
mem[127] = 144'h0f77f39e0e42f9510a2d00d903f8f2d9f413;
mem[128] = 144'hf1e1f65dffe9ffcffda6f753f1700187fccb;
mem[129] = 144'hf3cc0b8107b90d8cf5b2f28c00c1fc970617;
mem[130] = 144'h019ef11cf77df33001990dcffa0707cd0553;
mem[131] = 144'hfaad08e0f1c70574faddf88c0220f1430edd;
mem[132] = 144'hf5fbfc5ff7c2f37905c7f17105f4f76d0ec2;
mem[133] = 144'h04a6f9610d9cfab2073b0f72fe7b0c20fe5a;
mem[134] = 144'h0c6108910cca0fd302e4f9fef7f4f4eb0ec4;
mem[135] = 144'h04edf50e040bfb03f8a40ecf0372f52e0414;
mem[136] = 144'h0db1f95aff920a2c03fef632fe0cf55cf0c5;
mem[137] = 144'hf42dfba0f6a00479f2e2f681fa33f143f892;
mem[138] = 144'h0a200066068e06a8fe92fbb70be8095cf9a5;
mem[139] = 144'hfde8fbab060902040e5df6a8fa63069c0dd5;
mem[140] = 144'hf5abf7acf363fbecf67ff6170cde05450be3;
mem[141] = 144'h0584004603e0fa3f081805d50806f4b20c7e;
mem[142] = 144'hfe48f6ecf5b4f24cfebe01ba05fbf59afa96;
mem[143] = 144'hf3e80984f1dcfd44f983f4edf3550cabfb3a;
mem[144] = 144'h04c30ac707b9fcaffcbd01b8f38a0ae8f04a;
mem[145] = 144'h07d1f824f4fafe6d021f0b30f8daf038fdb9;
mem[146] = 144'hf3cffcb3044b09c9f828f2fc036f0ab8074d;
mem[147] = 144'h01d1faecf30af6bb05370d98019ffde90236;
mem[148] = 144'hfc75f214095c04340d970611047a098afcf9;
mem[149] = 144'hfc54f1bcfc2f09c1f48a04c7f8abfc080442;
mem[150] = 144'hf352fc97f9690410071ef99a08ee06faf254;
mem[151] = 144'hf1e1fcd200c60a84fb54f3660aff02330b25;
mem[152] = 144'h0b060ed309e90c6af0c4f2f1055709e6fa91;
mem[153] = 144'hf33707330922fb5cfbe3095a0bda0d8ff871;
mem[154] = 144'hf8adfb2efd9608e4f5bf0345f8f9fc7d0267;
mem[155] = 144'h0b310ab3f347f26801def5c3fd5af8b908c1;
mem[156] = 144'h0a0afddaff3a0f7f0c67fe2ff3fc0be8f5cc;
mem[157] = 144'hfda90e620beafdf60253f488fb1ff8a20862;
mem[158] = 144'hff050cec08aaf30000fff84308f6ff54f098;
mem[159] = 144'h019d096608530d0df07ffa15081cf41ef56a;
mem[160] = 144'h08d808c9f05e02ff0957f1480c32f30f0c3b;
mem[161] = 144'h02240c6ef90808dcfb530d3bf2c3059bf497;
mem[162] = 144'h02b10f43f357051af261076efbf906e9f8f3;
mem[163] = 144'h0af8ff23f7a3fefe006402c3fab9f58f027b;
mem[164] = 144'h0c52fdd50991f40bf955f98af50bf79c05ed;
mem[165] = 144'h064f0632fbbcf483fd62fbf30a690a52f6c0;
mem[166] = 144'h0dc7043d0a02f2880cdefeb503390336fc12;
mem[167] = 144'hf5930669fcb9f478f17e09bef0f306310cce;
mem[168] = 144'hf616fb690fc905c3fa87fe330db204aff98a;
mem[169] = 144'hf71c0b27f00a01dafb2a0678f46ffa0ef665;
mem[170] = 144'h099cf80ef45df810f01b0e96ffb4ff0bffab;
mem[171] = 144'h056e0c960e29005dfede0867f4f9080e0f27;
mem[172] = 144'hf81e0be0f63c06fa0714fb7d078a06ab029a;
mem[173] = 144'hf3010a7a01e3fabf058104580eca0ab705e3;
mem[174] = 144'hf958f2e50e8a0bf4f863fffe0398f6bd0cc0;
mem[175] = 144'h0e99f3c1f7180c320edf06270d66ff6d0f52;
mem[176] = 144'hf2c10cba0cd90482fb1700e80f4cf1f20e4a;
mem[177] = 144'h0d8cf48909d8f7a20cf8f580ff02f0680d77;
mem[178] = 144'h03de0121036efe6002c3f1be0d8b0c4302d2;
mem[179] = 144'h040af30308f5f18a097601290f99027a0dfd;
mem[180] = 144'h030c0612f68a0287ff350fbdf9450255fcf8;
mem[181] = 144'hf2260c61fa510158f6b50748f1a0f4ab01ec;
mem[182] = 144'hfbec020f021cfe33f3fe0a33f649006302db;
mem[183] = 144'hfbe5fcfa05d8f2b9fe16fe90fdc905f0f3a6;
mem[184] = 144'h09a8f598fd190cce0d24f97e04b400fe069d;
mem[185] = 144'h013505260ad5f6a9fccff2610e1ef169fa21;
mem[186] = 144'hfdfd0a6100cbf9c20d0c0faef374f51cfcc7;
mem[187] = 144'hf2500508f930042bf636f2f4f0be0121f288;
mem[188] = 144'hefe007f405b50f73071603e40ed4fc9ef1dc;
mem[189] = 144'hfbc9fece0049f31ff700f5c00df3f70d0d6f;
mem[190] = 144'hfd2a0cd4fe39072ffdaffed9f550012ff777;
mem[191] = 144'hf505f915f5fa0963fe38f8590443f5de0dee;
mem[192] = 144'hfc76f32b033cfe9bfc8ef7580ca407720ee5;
mem[193] = 144'h0791f4fb0fbdf98a0a060c8301e0f327effa;
mem[194] = 144'h07ca0d180c59010e058e082df1c8f524fbca;
mem[195] = 144'h032af1e80bc8ffd702670deff4b3f617f1f6;
mem[196] = 144'h041a0035ffbcf5e3fc86f5e2f65a03d20fd6;
mem[197] = 144'h0d9a07090cbf0bccf8fb0d5f01b00326f34b;
mem[198] = 144'hf511fb3a0ddbf9be0843fe57fc000aeaf6e8;
mem[199] = 144'h00090807fd7c0cf801dd03df0c6c0ba6f279;
mem[200] = 144'hf8a302d0f1a10b9bf2b5012ef53b0c62fd22;
mem[201] = 144'h0be9047e0a1f0eb8fed90bb002a5f781f0a4;
mem[202] = 144'hfd62f8910d380a200503f221052101b9f00c;
mem[203] = 144'h0faa08c5f97c0f5e078afc1f06c7f3c70303;
mem[204] = 144'h04c9fc220e6b038a03d9f219f1cbf45805d3;
mem[205] = 144'hf2f00575fca9f3b0fc3efb8c0bedf112f729;
mem[206] = 144'hf05702cc0463fe89028bf5200734f32af5ff;
mem[207] = 144'hf881019604d8f613f55ef2c1f4b40604f9ee;
mem[208] = 144'h041c0c0901befe98f290f6bf031efa70f903;
mem[209] = 144'h0749fe41f7050dc1004900a700e50c2209b9;
mem[210] = 144'hf9bbfa4aff8700d302bdfeb40faff6580969;
mem[211] = 144'hf6b10b8603f2f88cf207f80c0b2efc410514;
mem[212] = 144'h0ebd06f00b2cffcbfa2501b20dcffe7f0ac7;
mem[213] = 144'hf7eb029bfedf0e2105ddffc602f60ac4f953;
mem[214] = 144'hf069f6d3097ffe3ef2b60e88f1faf90c0594;
mem[215] = 144'h0c7a0b53f7750cd10ed908f7f97ff0e80152;
mem[216] = 144'h045fff8a0c8a04b7018403b9f78cf1a60d34;
mem[217] = 144'hfa7c029a06590205f455fd2504bdf23ef6cd;
mem[218] = 144'h0760086ef36cf44dfbcef74d0236f18ffa5b;
mem[219] = 144'h0898eff2fff5f45505500e52007df41a04e9;
mem[220] = 144'hf31906f30b09f73bf27401ea03c9001408dd;
mem[221] = 144'h0cfdfdb10453020b0c42f841f56e078ffe23;
mem[222] = 144'h0a55f9da0b36025708a90c9bf634fe66fd8c;
mem[223] = 144'hf7ebf7300c5c05e5f51cfce508cf07adf0dd;
mem[224] = 144'h0eba05180e020d2c09790c360c570524f8f8;
mem[225] = 144'hf146fb16ff60fed4fbb6f6a3f9f903470037;
mem[226] = 144'h0d54f94bfa0804260114f17005570c39f25a;
mem[227] = 144'hf820f244faa405e4f7f30d2e09300c3af32e;
mem[228] = 144'hf7acf9a30405fabbfcce02eb014d0824f7df;
mem[229] = 144'h05850e780043fea90868f5c9f9d2fa500168;
mem[230] = 144'hfbb90fe0f8daf8b705d8fe590f9900070558;
mem[231] = 144'hf91b0ad508c8f781f2e30d97faccf1ef0afd;
mem[232] = 144'h01c4f7e00cfbfce00b7cf96afc54f94f0465;
mem[233] = 144'hfbdbfa77087b0477fb8cf111f54e03490ee5;
mem[234] = 144'h0f14f2eef746065203cef8d1f49305cdfb8d;
mem[235] = 144'hf9f90bd70bbe01a000d80a76f888ffdc0328;
mem[236] = 144'h0427faeaf246f76ffd40f0720243fb440fc3;
mem[237] = 144'h0e8fff0f08e7000ff23ef7c8f928f70f0302;
mem[238] = 144'hf9cc002df642f1eef9c8f7ab035d0eef0d6e;
mem[239] = 144'hfa7407b007f2f5f20877f2a70bee05d60867;
mem[240] = 144'h0de202cb006c01acff4c0e900cf8f757f230;
mem[241] = 144'h09adf59d0afcf768feb60ba0f9dd0109f312;
mem[242] = 144'h09060bf3085e04b0ff1f0ae103bdfea00fb4;
mem[243] = 144'h04d10c3ff8ae07ef0d1101d200c6f00f037a;
mem[244] = 144'hfa2d0697f6dff69e0c15fff80e7b021bfd53;
mem[245] = 144'hf7d9fb520950f86afb5aff01fb85fcddf5c9;
mem[246] = 144'hfd8f06880ff3f7a30d0af2300085f36b0828;
mem[247] = 144'h024e056ff664003ff07b0d84ffc600a1f1bf;
mem[248] = 144'h01e80e01f3fb0115fd23fa6afa140232fe29;
mem[249] = 144'h08f5f744088af03af3c8fc3d049aff70f3a1;
mem[250] = 144'h0698065c0d270e13f52109bbf2530e0206a8;
mem[251] = 144'hf811f1fe0f3df5d6083c00b5fd09f09bf6f2;
mem[252] = 144'h09fff3980248fb7ef382f715f1690232fa9f;
mem[253] = 144'hf5220c98f50efcf6f9f50faf00780bb707c9;
mem[254] = 144'hf9090e080417f28ff44c05e60b9c071f0ad6;
mem[255] = 144'hf9a2f1dd0d3d0cd70408f660f492fe34f1ba;
mem[256] = 144'hf09004be0a1e0212f164fb410839f9aff4b4;
mem[257] = 144'h02a9f862f337f2960ad0f93b0013007d04bf;
mem[258] = 144'hf31508ba0e5df623fa4cf516f496f5c508b4;
mem[259] = 144'hfa7afc88f104fc760c5d0781f08905c209bd;
mem[260] = 144'hf9280d490f20f3560e7ffebff6f408e4fbd5;
mem[261] = 144'h0dfcf2b1f427f5e40312f22a0f94fd16f8d4;
mem[262] = 144'hfd6c00bd07400e81f4c8f5ec0e1bfa7d08f3;
mem[263] = 144'h0f8b0071fa800187f73e0f7df977fb700974;
mem[264] = 144'h0b3aff59f6a4f113fd00efd40245ffdffe84;
mem[265] = 144'hffcf02590a11ffd4fd7d0ccd0ec70c11f786;
mem[266] = 144'hff5a0b2bf0b6fc95f45e0f06ffe705030e18;
mem[267] = 144'h0dab0220f6cef1b6f7b8045bf526f6ee000a;
mem[268] = 144'h05a4f90ef8b7f2a9f467fd640abb072bf724;
mem[269] = 144'hfb5605b300d9f1e2f2730d240e8f0fc406ce;
mem[270] = 144'h01c20d9b0dbffd5a0bd001ecf68b001f080a;
mem[271] = 144'h0eb90366f143f40df67af0e3fe01fd160a18;
mem[272] = 144'hfa130b350499f964066ef2d20748f50e0748;
mem[273] = 144'h0557f53efe25fe45f3180d930961081a04ae;
mem[274] = 144'hf8d3fc97046b099afd91f37ef0e70701f002;
mem[275] = 144'h0081fe100bc601aa0f7005c3f83ef907f106;
mem[276] = 144'h0d600695012df4c0efebf4e004a1077d094c;
mem[277] = 144'hfa03ff49f6820625f5470d1b03bb027af76e;
mem[278] = 144'hf053fd14f92b0aaa0dd301c9f6ee04ff0391;
mem[279] = 144'h0dbe0e0ffad70433f1d00d2ef5ca00dcf05e;
mem[280] = 144'hf3210cf4012cf3aa04d4f2850f5907180c03;
mem[281] = 144'hf2db084b0317f9f8f51800490acdf672f71b;
mem[282] = 144'h0b65fcfa063ffbcef3fcefc200cbf39bf7f6;
mem[283] = 144'h025402a40fb308a00d3af329f795fb2b0f83;
mem[284] = 144'hf95af951ff90f534f3ea0906074afe440818;
mem[285] = 144'h027effe9f85cf23500820841083efd6704c9;
mem[286] = 144'h07bd0484f60b06370c550bf9ff2df493fc4b;
mem[287] = 144'hfc04fd840588006908b1f5a502030c81f5e3;
mem[288] = 144'hfe16f1e5fff4f47a0d7b079100bafe050873;
mem[289] = 144'hfbc3f72e02abfe44f64b0d810ddc06effb04;
mem[290] = 144'h0d080c3bff65f64a0879f899024b0c2b0c5a;
mem[291] = 144'hf3fafb30f7ec075dfa45f45d0fe70a4800b3;
mem[292] = 144'h09dff4420ab50bee033ef84609280ee4f107;
mem[293] = 144'h0dccf51df5f4f3f7f7e5004d0a06f418018f;
mem[294] = 144'hf9bbf6b202ed0c320e080e3c05f90c0e09ea;
mem[295] = 144'h014f07acfde602450006fdb00448064bf96b;
mem[296] = 144'h0bf1f421002b021bfa480e76f872fefbfc16;
mem[297] = 144'hfac8f686f280056dfa2b035500d8056504c6;
mem[298] = 144'hf6a60f5cf55bf1bc0e9bff0507fbf4dd02a6;
mem[299] = 144'hf2a10a1d0584073af96a062c0820f517f029;
mem[300] = 144'h068e0a45fc5b08b40c4ffb5e09a20f3d0ba4;
mem[301] = 144'hf751f0fc086df425fcef049d00bff7b002b2;
mem[302] = 144'h0e65f2c3f4a7fbb20d6cfac40bb4fbf6fe0f;
mem[303] = 144'h077f05de0dd2049103250b82faf401a1fc14;
mem[304] = 144'h0b2c017b08a6fa45fedef12b0678057e0ef3;
mem[305] = 144'hfc8503550ce00c30fc0efc2cf58f0be5009e;
mem[306] = 144'hf37cfd73fe06fcff0fd7f9e1f0cc097e0b91;
mem[307] = 144'hfe7cf0e30f8603620f8b0f1d06bbf93df986;
mem[308] = 144'h0f47054b0a19070a091f070efcce086a097c;
mem[309] = 144'hf861f831efd5f4cff19ef80b0308f32d01c5;
mem[310] = 144'hf8a609c107f00da1fdcf0395fecd0858f948;
mem[311] = 144'h076407320abf00ecf74308ba04a8fac7f6ce;
mem[312] = 144'h073ff9e201670f9ff4aaf5dc02700da50665;
mem[313] = 144'hf1d207da0055f3e0f80a06b000f60eb30df0;
mem[314] = 144'h06bf022a027ef40d0372ff2607a2f9470852;
mem[315] = 144'h0d4203acf904068d0c25f9350acd083cff1b;
mem[316] = 144'h0526fff90d4bfe75f5d3f6ac01f308c707cd;
mem[317] = 144'h09abfb180bf90a64f8200fa104f9f22d0dc8;
mem[318] = 144'h096a0e23f4e8fdd4fbb2f2a8f782f1f70733;
mem[319] = 144'hf2260c1a0e1c08dff5fd0afa075002d1fe5b;
mem[320] = 144'h0aed0e2404d70376050efb8df9acf02505c7;
mem[321] = 144'hf4a4f0b306db0ef2f85ef1280e4bf831f871;
mem[322] = 144'h0909feaef5bcf788f868035706880ac1062c;
mem[323] = 144'h0f8a0729f3ff02960396fd5af6c1fc76051d;
mem[324] = 144'hf584fc0401b9f013044b0fa60a8b021cf108;
mem[325] = 144'h0ab7efe00b5f0673f54efcedf1b5f47b03c0;
mem[326] = 144'h0b8efcbafe2f0e46f7bb09cdf7f309bef819;
mem[327] = 144'h0cb7f3c2097e0d660f80fd3bf0b30f0a0f57;
mem[328] = 144'hfde4fd10f08efb78fe280634f92d0e67f4f7;
mem[329] = 144'hfaeefec600dbf06cf842fc5efec50aca0c12;
mem[330] = 144'hfabbfc6e0b96f339fa3af3fbf57d0d760eb8;
mem[331] = 144'h050f00f30d94f8030a9cfcb9ff180a5f030d;
mem[332] = 144'h0d1600f4050afdd5f92e03190caef650ffdc;
mem[333] = 144'hfc0afbd701b2f22ef03df2cffbf1fd920446;
mem[334] = 144'hf3b1f9a301a3f9f4fae3076b0dc70495f85f;
mem[335] = 144'h0abf0fa5f3b208460199f4a0078dffae00e3;
mem[336] = 144'h035a0611fd6407010c55f64b04c20bf9fc13;
mem[337] = 144'h0f0b02320eb3fb64f12b035df5e30f210ebf;
mem[338] = 144'hf33bfd7efe2cf8b5095805a2f6d201160c4e;
mem[339] = 144'hfcc6fb3e010df24204ddf25904850e6b0320;
mem[340] = 144'h09c40014fdb609eef3be01bef5370330f097;
mem[341] = 144'h04ad0845f04efcd509680ea6f1d2fe07f005;
mem[342] = 144'h06d7f34af14df1fbf24501ff0aadff4ef1ea;
mem[343] = 144'h0da802c3054df082035f052802aa04b4f2f7;
mem[344] = 144'hf678fced08320d750f3d05710d4205690d68;
mem[345] = 144'h06690f79014d010600d0f94907f402dbf406;
mem[346] = 144'hf4cd05c30a9f0834f927fba3f97909c807b8;
mem[347] = 144'hfeb5010cf0f6000b0053f15cf917f346ff87;
mem[348] = 144'h0ca3006dfd73f080fedbfdc201a1fa020271;
mem[349] = 144'h0c9df8eaf929f658fed6f52a01fefa36f725;
mem[350] = 144'h00bdfafa0da3f3640d77f028fae60005007f;
mem[351] = 144'h094df3f3f2baf0f4feef0405fed2faf9079e;
mem[352] = 144'hf447f200fa350c9bf59bf016fb2bf308fded;
mem[353] = 144'hf270f78a08940f73fe330312ffcf0585f334;
mem[354] = 144'h0892fe91ff9ef045f44e0f6ff828f6b2febe;
mem[355] = 144'hf1fb0483fc1dfbea033df374f3de0abaf1f8;
mem[356] = 144'hfba9fcc4f95af7d906bc0499f68102ebfe51;
mem[357] = 144'h044d085ef018f7f9f1f104e6fdb3feebf601;
mem[358] = 144'hf7290bcc0e950d0c0b4a0136f952f91d071a;
mem[359] = 144'hf8faf6eff808f694ff3df64105150e2606f5;
mem[360] = 144'hf4f80ee8fe17feee0abefc4bf3a4004cf4b0;
mem[361] = 144'h04b7fc4bfbfefdb2076a0fa20d9f031df20d;
mem[362] = 144'h0669f65cfbec0bb4f325ff79f924023ff025;
mem[363] = 144'h00420f25f2f2fd0ffa5ff76f0836faea0d12;
mem[364] = 144'hfa57f5c10e44fcb609f50824044ff6a2f953;
mem[365] = 144'hf4a4fd17fc33fe67f49c08f30c34fa0bf559;
mem[366] = 144'h0e1ffd36f4f604b00fe8faccf28ef542f160;
mem[367] = 144'hfae90441f218f4c50981fe18f6520791ff71;
mem[368] = 144'hf79afa5d0ca9f9d10983059f0499fc8afba4;
mem[369] = 144'hf8bffd65f257f2af04d2f3f9ffabf101f3e8;
mem[370] = 144'h052506400b8e0daff1230fb20eac00f8fbcb;
mem[371] = 144'hf95108b00913f10909860f1c01c40c7c0c84;
mem[372] = 144'h01fa0ebb09af0c50f32005c9fb000ec50acc;
mem[373] = 144'hf98af07e0ad1f96bf303089e05fd05edff21;
mem[374] = 144'hfa060388ff750bcb0307f049f3b1fe73fe46;
mem[375] = 144'h078ff119fb2902a50980f58ef243046609bc;
mem[376] = 144'h0754f5e3fb34fe73f893089fff2d0993fa84;
mem[377] = 144'hf4960f84096505ccf3400ca00cc3ffb8f136;
mem[378] = 144'h0d91f5d103dd0fe1067d09b7091d01e9f8cb;
mem[379] = 144'h09b6f432f5480b62fe800780077af034f736;
mem[380] = 144'hfaa7058f09fe063afa5b002afeac0b88006d;
mem[381] = 144'h0485f6b4feae0fa1f720fbc000090300fc7d;
mem[382] = 144'h0449fccef5a109850eb1fe020b4bfcdcfada;
mem[383] = 144'h03380eb4fb58f15af40905bc03640b3ff32e;
mem[384] = 144'h0aee0b13f4b90d1501b9f287f66b05b8fb3d;
mem[385] = 144'hf59f046d0114f2af0d730ddc0cd807f40609;
mem[386] = 144'h08bcf31206e10074fe850806f5cf0af8f277;
mem[387] = 144'h01a905a00d36fcc6035f024009350dd70e81;
mem[388] = 144'hf93af3b30fa30aaa02aa0e7df7f8fe210978;
mem[389] = 144'h04fcf3d9086f0101fdcaf3990584fb7cf08d;
mem[390] = 144'h0f5203c9f2a9f0590253f93dfc3df931f3f6;
mem[391] = 144'hfcae0ffafe630794fb980e8b0c4bf1b2face;
mem[392] = 144'hf99e082f0c260e90f877f8290991f6f9faa4;
mem[393] = 144'hf0c700a1fafd0f2d07a4f398fb40052dfb07;
mem[394] = 144'h090209f6f949f30c0b7705baf7a9018ff3c7;
mem[395] = 144'h07090240009807450be906f4f21103c9fa2a;
mem[396] = 144'h0890017f0a9c08f508ca0ab9f6cc0906f157;
mem[397] = 144'h017ef3fdf5160548f0eff235ff040496fe8b;
mem[398] = 144'h0aa70c310c130357f321f55b095607c9f5c4;
mem[399] = 144'h0f140a29f3570fbdf28c0764023ff313f89d;
mem[400] = 144'h07a7fe4901f201a408f6faa902c0f4baf5cc;
mem[401] = 144'hfff7f2680b450e5cfa66f1d009ea0a05fb1a;
mem[402] = 144'h0db80742039ffed401d3f8b30959f6d90fdb;
mem[403] = 144'h07a6ff84fb8b04f4fbf0ff65fd36f413f5c6;
mem[404] = 144'h06fd01f5003ffb560b08fb89fb0f06200df1;
mem[405] = 144'h0f0cf27d0b4ff537f053f84cfb58f9d4ff28;
mem[406] = 144'h0e1cf97bf1a8f7a0fb0d04bef69dfb530694;
mem[407] = 144'h08dcfbdf066100af04a10f3e067efd8e0eb1;
mem[408] = 144'h01f60e300e81040200d6f68a0a530c430d50;
mem[409] = 144'hf5d206d2004dfabd02df0c670b26fc4407e6;
mem[410] = 144'h0c850614ff37f579f045f09001780e0af430;
mem[411] = 144'h03ecfd950199fb1afa3705df0f9af6d6f19c;
mem[412] = 144'h0c88f51bf04705ec0130f0ad0fd3f6f0fc83;
mem[413] = 144'h07a5fbc50387fe5a0e07fc6dfeaef1020af1;
mem[414] = 144'hfcb4fa8ff372f06dfbebfe5c0275fcfe0976;
mem[415] = 144'h0cd20c59f80ff53af5720ae3029103e30b93;
mem[416] = 144'h0f5ef2a2fe2af3cf0f03f868fe4d08e50a89;
mem[417] = 144'hf42aeffa013106870474032706f70c1cf067;
mem[418] = 144'hf5a9f429f2df00c0f7630e87f14806ef0bd5;
mem[419] = 144'hfa3009fc0d270268f59604a3f2adfb25f25a;
mem[420] = 144'hfa83fef3f61bfa16f762ff030f90f78cf671;
mem[421] = 144'h0671f27f0ddef09cf58009f5ffb8f151f273;
mem[422] = 144'h08bc05e204300dc20bab0be50046039e0f6b;
mem[423] = 144'hf0ae0eb6fff80ea6f2520e1f004fff210933;
mem[424] = 144'h01c5023202900b5a062f0937fbf706fbf7c1;
mem[425] = 144'h0010f847f9d7fc42f832044907e9f8390e8f;
mem[426] = 144'hfb61f29e008eff8105a0f444f6f90512fc32;
mem[427] = 144'h0c00f2490fba03d0f5e0fadaf145f42b0216;
mem[428] = 144'h05a3f1f000640ca80b6408f1f845f9550ba5;
mem[429] = 144'h0ad20d12fd52f206faaff156093806010110;
mem[430] = 144'hfb3f00e400dffd5b039f0978f5170a790bde;
mem[431] = 144'hf7f9fcfe0d15f105f99109e6f109088dffd1;
mem[432] = 144'h04b302e10688f176f3f1095efa1df3ef0a88;
mem[433] = 144'h078af62cf22a05790690fdbf0275f244f77a;
mem[434] = 144'hf09bffabf37cfac5f486fcfcf9d10b64eff4;
mem[435] = 144'hffbbf258f3cb0f2cf1d6f6de02bc06d10f9d;
mem[436] = 144'h05a9f516014af4e6f63af41403f708a80b93;
mem[437] = 144'hfb1e02b2f074f0000f3a080ef5530e3cf805;
mem[438] = 144'h0a61fd97f9affe9bf20706b20097fd43fdf6;
mem[439] = 144'hf27ffd56fb230f70f3d0f98109f50e6bfed1;
mem[440] = 144'h0698f267005efaa0fd420b4ef9210a50089a;
mem[441] = 144'hf6730ea20ff107c7f21a0e2cf70b0051fcda;
mem[442] = 144'hf0f80503f5080de2f5460434050ffa3e0706;
mem[443] = 144'h0433f91cfc63f99b05aeffbe08ae0b7f0b28;
mem[444] = 144'hf97bf44bf104fcd00da9fa60f6f90be409fe;
mem[445] = 144'h0e3708e709ba04080b590b1cfea3fcddf229;
mem[446] = 144'hf670f468fd950ef5083af2c007560dbd0d5d;
mem[447] = 144'hf720fbe1f47d018406d3fd2ef5c3ff940938;
mem[448] = 144'hf494fec10df5f155f2b1f6f9058ef943fb36;
mem[449] = 144'hf89ffb03f048ff360f5d0996fcd405d40476;
mem[450] = 144'h0a72f8170233faa105a5f6e90ec7fee205c2;
mem[451] = 144'h040cf0e4f11dfe1cf4c5061504710400fdb1;
mem[452] = 144'h0aac00cef7f5fc6df135f28d0314f51ef82f;
mem[453] = 144'h0774ffa4f60f00030160fd83f38ff2630299;
mem[454] = 144'hf1c0076307acfe2ff65907430d610d79f568;
mem[455] = 144'hf788f50909cd0976f5920d6bf1950220fd32;
mem[456] = 144'h0f58f1bffa10016c0347f95efbc2f37ef3f1;
mem[457] = 144'h0a850d71015706e5039ffd9a0ac7ff220668;
mem[458] = 144'h0b2e001cff8f00320223fd10088cf1200262;
mem[459] = 144'hf9410d28fa4f04820b8df7c90ee9f5e507ec;
mem[460] = 144'hf0e00ebafe83ff6efaf4ff2c0da2fb1404ac;
mem[461] = 144'hf7a0fcaa0304f5c3efd1f97efcfd03aefb24;
mem[462] = 144'h0e3b0d96f500fac5041ffd41042f0119f854;
mem[463] = 144'h087901400a26fa380211f432020ffe62f924;
mem[464] = 144'h0905ff260e61f1340282074df53f04dcf169;
mem[465] = 144'hf6c40a76025ff44b002a0831fe4afe1d077f;
mem[466] = 144'hfef902d9feae0f8afb5303fcf85cfeab04bf;
mem[467] = 144'h080ffdbb0cda08c4fc11f7c9f3ec0a940849;
mem[468] = 144'hf15cfa3bfc87f9ac0a6901660279f284f1e8;
mem[469] = 144'hf950ff9605fb0d540d3d060102430e36f4be;
mem[470] = 144'hf484040f0203f2410ce008050e3efa43f040;
mem[471] = 144'hf8daf847f54f0737f96700cbf85ef0f9f01e;
mem[472] = 144'hff5e03f4fa2603eb03200a380f6d01ce0495;
mem[473] = 144'h0561f519ffe30f6bf230fda7f7210ea2003a;
mem[474] = 144'hfacbf5410ab5f6dd0819f2420e680ee80d1d;
mem[475] = 144'hf55ef32af4aefb240109026ffd28f333ff37;
mem[476] = 144'hf5460183fc040d24013406aefa590db7f79d;
mem[477] = 144'h0777f807048af1e4f84702d50ad3f9000d76;
mem[478] = 144'h0b51074ffc48fe7c0d25025a0937fdb30f0c;
mem[479] = 144'h0f8c02c904980c08f7acf42bf4c5f7d30d7f;
mem[480] = 144'hfd050004f81bf8d90c1802b906610dec00ea;
mem[481] = 144'hfd91fc9001b80752f92a0bd3fe3ef5bcf1fb;
mem[482] = 144'hf33df73b0163ff1a0051f072f3da0e21fd01;
mem[483] = 144'h060af4920d9b0214f042043b0b8df7090d87;
mem[484] = 144'h0eda0900f69a0a21f0ca0582fce4f9ee0efa;
mem[485] = 144'hfee804900f0a0e350f2005fcfbe1f76bfd0b;
mem[486] = 144'h001d0d3106c8fff3f620f1f70e6407d4f8d6;
mem[487] = 144'hf8d3f9d3f6ddf4d00a1e0b5df7970985fc01;
mem[488] = 144'h07b9f628f23409fa0afcffedfdce0bc7fb98;
mem[489] = 144'hf06cf234f223fdbdf3e40c370802f2950017;
mem[490] = 144'h0783f1710508f174f4fd0ba6094cfebb053b;
mem[491] = 144'hfbc003a3f4c0f287f188f6f6f9e7ffa4fee3;
mem[492] = 144'h0ece02f003f502190b7909c20c0e099e0fa5;
mem[493] = 144'hf84ef0e70d5a086df0e6f90cfc31fb31fd07;
mem[494] = 144'hfe090b66f866f3b9f1050cf1047af641f44e;
mem[495] = 144'h00360d33f9cff62ffd6001cf07a40b630869;
mem[496] = 144'hfd1ef628f80a0e5dfde309e60ceb050f0fac;
mem[497] = 144'hf7dd019e006af03bf5d20e3d071b04affae6;
mem[498] = 144'hf2b80e84f13407de063bf14d035f0401ff3d;
mem[499] = 144'hf45c09cc02e0f0920edc0e9dff9afa360be8;
mem[500] = 144'hf43af2030925f8e9fbbf0afa0174fa60f218;
mem[501] = 144'h08300ad20264faf4f3e8f5d8fb6ef2b40c92;
mem[502] = 144'h0586f880049efc1cf42608e2ffd7f690fe46;
mem[503] = 144'hfa64f62f0b0d0b0f05def8a90935fac1f16f;
mem[504] = 144'h00f20809fde7fd99f897faa609fb0a200ecb;
mem[505] = 144'hff57f67bfdf901a009700c26fcc8f684f2f9;
mem[506] = 144'hfe8dfca9fca704b1ffd7fb3dfb3402dffdf2;
mem[507] = 144'hfc50febdfb7400f7f01a01c103340752f8d7;
mem[508] = 144'hfdaafff6feb706def2c90d47fa4f0b62ffce;
mem[509] = 144'hf5890bee06dbf6a70907f9c70c0a044afbca;
mem[510] = 144'hf5c50f69f855f15a0b45f0520a5602e4f470;
mem[511] = 144'h02a2fa150be4f9510894f1870017f41900fb;
mem[512] = 144'hf773fed1fa73004702ccfb8bff370534f34b;
mem[513] = 144'hfc66f316fbe60aa10913f4c6f520fa020c4f;
mem[514] = 144'hf387f1c50284054202edf5b6047d0993fc5e;
mem[515] = 144'h0cf7efd4f1b4004efa24070bf8c8f6ee0ed1;
mem[516] = 144'hf46103eaff1b0b1ef58b02f308def5a4f74e;
mem[517] = 144'h011af05901d50130f005f042f2d9072b0b55;
mem[518] = 144'hf575f03ff9a0faf908bef0570238f9a0f121;
mem[519] = 144'h05fef3adfdcbf1700e2f0dfaf5f3f9d60ad6;
mem[520] = 144'h0f68fa6202cef148fc21f48cf1d9f228fc0f;
mem[521] = 144'hf3810147f5700ca7ff5bffc6fac3f5cc0316;
mem[522] = 144'hf481f23cf424fcb1f2270b8e047206ed0f91;
mem[523] = 144'h01da0ec70694047bf741f840f41a0bb30212;
mem[524] = 144'h08f3fa72f73a0459f20df006fe2500c4044a;
mem[525] = 144'hfe24044c07360573012801e80789ffc80b10;
mem[526] = 144'h0273f43bf5ea0fe4f03e0876f108fe47fee7;
mem[527] = 144'h0b23f9c5f95b037809610779f4450fee05c9;
mem[528] = 144'hfe04048801240a1a0d2af465effc067a0a97;
mem[529] = 144'h046af463033a0c51fdd5fc0f0976f6a60071;
mem[530] = 144'hf544f5d2040509720031f6680bf8fcd5fe5e;
mem[531] = 144'hfc17f3130c2dfd070e8e0ef7f9e5f0e0f97d;
mem[532] = 144'h04e00462ff22f63c001ff1ffff0df7dff10e;
mem[533] = 144'h09cc0aee0df9fb2cf073f0e70f83081c014d;
mem[534] = 144'hfc7907430165f02f06d2fb270faef890f1d3;
mem[535] = 144'hf9f50e230e0a0497075f00990b35008ff1de;
mem[536] = 144'hf3c6fe83faf9095b0b6ef862fda4016402c7;
mem[537] = 144'hf538fee2f151f3b4f1baf9fef4ac0a51f034;
mem[538] = 144'h08c50290fcabf70df3f1fa99f1f5f055f76b;
mem[539] = 144'h03bd0f86f6fffbdbf6b6f143f5cffba60978;
mem[540] = 144'hfe0f0ee9f95202e40fc50862000dfa1c0ab1;
mem[541] = 144'h07700df7f82708b6fbc1f70107f101ed0961;
mem[542] = 144'hff4c0bfffd18026ff165043e08d2f2920418;
mem[543] = 144'h009b0371f825f50f0090ffcdf6880092f457;
mem[544] = 144'hfafe0a87fa960946f54d05fcfab903e20c18;
mem[545] = 144'h009c0daaf18ff498f1c90f9c08df043bfa53;
mem[546] = 144'h0f0403c7ff44f8b808d406d70c9efa0ff0b6;
mem[547] = 144'h00c8fd790b2af708f0ec0847053805c106b6;
mem[548] = 144'hfa8cf29806fbfb5cffdf078ff2ce0fbdf417;
mem[549] = 144'hf4a4087b05da00190f13f319fd4f0c6afeb0;
mem[550] = 144'h0d2809be097d0882fee1053402020623f15b;
mem[551] = 144'h0c83fddf0907fe23f143ff4c0fbf0265f586;
mem[552] = 144'h0e3efe86ffe60913f69b04b4f06b0f67fd99;
mem[553] = 144'hf508f8e8f5f3f2770548fac1f7e5f98b0c8f;
mem[554] = 144'hf9e6f272f6b4f18504ff061af2e50a59f72d;
mem[555] = 144'h05960a64f45a0313f85df270fe560231005d;
mem[556] = 144'h06c905600c230797043e026e010f0a8ff745;
mem[557] = 144'h0bf90876f4b00836f15e054000aa0738fb13;
mem[558] = 144'hfc720cf70869fd5bf66308300a8bfb68fb82;
mem[559] = 144'hf1190876033001e300e5faba0d9405e80b1f;
mem[560] = 144'h05ba00520c0604b00d95fec4fb02f4c9095b;
mem[561] = 144'h09b00520003df3580d38fa6f0587f128007e;
mem[562] = 144'hf926f953f523f91505edfe2bf1b3fc1ffd9b;
mem[563] = 144'h0fa2f7860233f75ffcb500cd0000f9280cd5;
mem[564] = 144'h0f480b15f418fb120badf4ea0de2038f05c2;
mem[565] = 144'hf66df940fa98f2ddfb860afa087f034bf4c7;
mem[566] = 144'h0ecbfc0d05b20f10fb6e02a403a6f55604f8;
mem[567] = 144'h03880fe70a7ff06d0e3df89e01f504820fa4;
mem[568] = 144'hf43cfab3fd2205bbf466f285fc35093ff0f1;
mem[569] = 144'hfb4c0d06fcac0af6f1b9ffd209f101d1f1cd;
mem[570] = 144'hf37e0623fa26feedff8504a605fa0413fd66;
mem[571] = 144'hfc96fff207e0fdfef38a0abefa66f8010fdb;
mem[572] = 144'hf523f389f6ed08ff08f7fa75005af0410ad8;
mem[573] = 144'hf27b063df0190d290050035dffa5fb3508d8;
mem[574] = 144'h0069f942063609960a7e0701fb73f8550de8;
mem[575] = 144'h0ccaf6f303e7faadf9c8f5bcf1820267fb56;
mem[576] = 144'hf4cd02eb02baf506021c00fe04a707940971;
mem[577] = 144'h0921f24bfb34f0e7f34d00a0fdc10b15f5d3;
mem[578] = 144'h02f0f42f081f06e3fa070ad7081306d7f362;
mem[579] = 144'h0ea90e9afebdfe07f8d1fe34fe35f0fb0bf9;
mem[580] = 144'h053a0b940e6c02b8021af2a4f165ff74f0e7;
mem[581] = 144'h08450650fae0f8d8fe18f31a07a3ff49ffa3;
mem[582] = 144'h082cfa230ef9fb83f41c092df49b00d9f0d1;
mem[583] = 144'hf65cfd33f8cff4bc0e0903bdfbb901a9faf1;
mem[584] = 144'hf3b00628f8e60e680b9909befd13f78df88d;
mem[585] = 144'hfe2bfae5f4f8fa500963f48ef88c0c79f604;
mem[586] = 144'h0f4cf36a0aa80231ffb701c40d2e0fd2f63c;
mem[587] = 144'h0ce50b150d9ef5dcf77ffbe8ff160c2105b4;
mem[588] = 144'h041606ca009bf6bcfac1f9e1f1ed0822f3f7;
mem[589] = 144'h0230f2e902980cb70ca4092af45f05acf173;
mem[590] = 144'h037e0201f6cefb81fbca05b5f4d8fc69064c;
mem[591] = 144'h01b4fe7209eff4a807a80494fbd6f9f907ae;
mem[592] = 144'hfcae0307f9d3fd1102cd01ad0c2e06b5fd79;
mem[593] = 144'h0d3f0c73f4a0f7370503f3a2fbb4037b0547;
mem[594] = 144'h0b31f5e80966f5d00a94fc750b73f62ff150;
mem[595] = 144'h0a2afbd4f2250d6efb8c046dfa6af9010a83;
mem[596] = 144'h0d4c08470783fe94f56ef18b04c2f7d10b42;
mem[597] = 144'hf99d0d380daefc17fdb8fa250b8ffa34022d;
mem[598] = 144'hf2570c8f051ffde9f387f275f9cef66f0b8c;
mem[599] = 144'h0e410076fc4503c9f2e20e820fdef0bc00dd;
mem[600] = 144'h0d2a040c0ac7fc9e08c702ad01eefc70fafb;
mem[601] = 144'h0ac90150055bfeeb03e7f13af56a0c06f74f;
mem[602] = 144'hfa4bf28f01240759fb7e0daffcdff1b5f45e;
mem[603] = 144'h026f0c2f0fa2fb72fcb0ff8ef180f15efd8a;
mem[604] = 144'hf2420ca40cc70ec2ffef05d60347fb5f05a8;
mem[605] = 144'hfa2607c8017d02c1025df1880ef40f2c02b4;
mem[606] = 144'h0510fec4f2b40246fed1ffd2f0ee001e0642;
mem[607] = 144'hf0ab0b36f27305dcf82c02a7f0e2fddef764;
mem[608] = 144'hf0380837fade069106f50401f8d308510447;
mem[609] = 144'hf90e0a3b03910ba3f72009270d1b0028f195;
mem[610] = 144'hf7d40e83f9160a9005110a91ff69ff70018f;
mem[611] = 144'hfd54ff97fc16f9f908d9f9a901e4f39cf11e;
mem[612] = 144'hf49d0e0103cbf1020d0ef29107740f2af907;
mem[613] = 144'hffa00df5f99e08e1f65d073609b9fe9afae8;
mem[614] = 144'hfd4dfec7f7e20ba2ff4af26b0737f505f640;
mem[615] = 144'h025cf49b0da70da3f422fde80430fdc00df8;
mem[616] = 144'h0e33f37cf179f3d8083007ca0c06f3db0a87;
mem[617] = 144'h0d31f224f58d0692fd3c0c3a0f20fce9f1e2;
mem[618] = 144'h0f5e0e04f4e30ed1f48702a1f585fa14f831;
mem[619] = 144'h0291ffe702230d6808af0bfef08e02ea01af;
mem[620] = 144'hffec0f490b2bf6f2fc6bf480036c02b10ee3;
mem[621] = 144'h095df2f7fbb0fe18efdaf3aa0c1ff9b1f4d5;
mem[622] = 144'hf9fd0dc8fd4a0e4af16107aff30209170b1e;
mem[623] = 144'h0dd40392f345f7130b680fb40181f0ccf4cb;
mem[624] = 144'h07d10745fc27fe160cce0c6d05b505d30eb6;
mem[625] = 144'h01da07310f6bf96f00420a9803b50a6df915;
mem[626] = 144'h0747f97f0013f55702b407bdf25ef3ab0365;
mem[627] = 144'h0a01f87307adf8f8fe23fe24f066f24a0cff;
mem[628] = 144'hf35404b901f8fc170528f6cff2fa06e4fd80;
mem[629] = 144'h0424f870f13af498fed7fb80007cfe71fd51;
mem[630] = 144'hf57b0d49fe65f2df0d7cfffa020d0838f763;
mem[631] = 144'hf49dfe6efe24046bfb9e0bf9fe59f6e5f138;
mem[632] = 144'h054df1d1077204dd02dc04b7ff66f336fc0f;
mem[633] = 144'h0876fe370bd6fe72f470f2b2059cf1edf4e3;
mem[634] = 144'hf60bff72f44100020639fcfdf1f70f54f92a;
mem[635] = 144'h0fc600f70483f48801760f10f2a4f799f7c1;
mem[636] = 144'h0b090aa80e2602510a6ffabdfc22ff81fc4b;
mem[637] = 144'hfbe0f98c0e880adff126032e0130f1480dfe;
mem[638] = 144'hffcbf0be0bbc025afa41089ef9b4fc8df87d;
mem[639] = 144'h05eeff3f0df206c30a1b06190c86092ff1fb;
mem[640] = 144'hfe7f036d0f6af80c0c41f2c2010cff4f0082;
mem[641] = 144'hfa28f678f6fb0bf7f4b3f693fb4007bf0a20;
mem[642] = 144'hfcabf78ff7600e7af06e0286f2d2f43f0791;
mem[643] = 144'hfdfd026b00adfb98f19e051f018902940417;
mem[644] = 144'h0e110fdff742016fffe2fc680921065804dc;
mem[645] = 144'hfd40f4b60229fc6b05e8001ef81f02d0f5a3;
mem[646] = 144'hf816055af7f30e79f715f577f4a50d43f2ca;
mem[647] = 144'hfa580e85f8580d4ff42f064707970600f591;
mem[648] = 144'h01d6fd990e660c59f9f00edf0837fa780dc8;
mem[649] = 144'hf0b105db0875f9e003a0f5baf1ae0aeafc45;
mem[650] = 144'hf966f0a60824fbc7f0340072f20608ddfd2c;
mem[651] = 144'h0f5af50001d80f92fedd099c074b0b3ffa7c;
mem[652] = 144'hefd20844f4dc0176fc220ed70128f2f0f04d;
mem[653] = 144'hf0d3f1ef03b50d99f94101e00d57fd66f6a5;
mem[654] = 144'h0d7a0ad6f232f230f2c5f6b90edd0ef9f64c;
mem[655] = 144'h0378f93f0486fc5f01fb07920d44f8d607c1;
mem[656] = 144'hfcdc0185fae4f15ef42d076af126fe2ef486;
mem[657] = 144'h020701ae009604d1f7a8065dfc7a0f8001a8;
mem[658] = 144'hf9d904e8f5f707030aa6f4f2f63a0e1df80a;
mem[659] = 144'hfc060093ffe2ffc2f1770a220dcff03f0251;
mem[660] = 144'h0780078f0c52f2000a4cf9020d89f5980d7a;
mem[661] = 144'hf5fffba604980da3fe25f82d0c18075d0aae;
mem[662] = 144'hfd1af3d6084d0090f2a8f2ba016bf6dd0d2d;
mem[663] = 144'hfb12f0950762077cffd9ff1ff7bd047df53b;
mem[664] = 144'hf4d70d9dfa2af4fa041d0f23054807a600ee;
mem[665] = 144'h0d70f1e1febff07d0a65052eff05f75af589;
mem[666] = 144'h0ee403cd041a07f6f5420bf80cc006dcf668;
mem[667] = 144'h01d204a00c8ef623f46b00a6098408ab0a92;
mem[668] = 144'h03d6f499fc4804a70d6cfb4dfd02f1530318;
mem[669] = 144'h0eaafa1306200cfa0cd6fb4a074dfa87fcd4;
mem[670] = 144'hf492f098f2d2f4f7fdda03700b69fb05f3cc;
mem[671] = 144'hf6aef5d1008ef99f06360cd5f48dfbee0ded;
mem[672] = 144'hfa81f874060a0e97f7af0c46f99707d4f878;
mem[673] = 144'h0a18f68308cc018df575fdf20878f1f9fb88;
mem[674] = 144'h04ebf02309e0f44bf3a500ec08e70430073d;
mem[675] = 144'h06a10f520a900a0800fcfa35ff6a0afd079f;
mem[676] = 144'hf0bef1d60072f6d2f934f4ca020eff0df95a;
mem[677] = 144'hf22ff72107a3f7f6fd5b02770b220ffa05a0;
mem[678] = 144'hf771fe9400b5fa7c0039f6ca0401f565f536;
mem[679] = 144'h024af00901c6fc1d06eafc7509fffd6a08de;
mem[680] = 144'h064af36a0bb3010407f4067009e0fd3106f6;
mem[681] = 144'h02500238fd74f02df383f9eef23df1cff12a;
mem[682] = 144'h0c92f7e1065ffdacf550fec2fda4078dfadd;
mem[683] = 144'h086ef670f0a7fc98f98d0af8f65ffc4208aa;
mem[684] = 144'hf20ef1b60ff30789fc880be2f044ff640506;
mem[685] = 144'h0d140a00fef0fc84f5fb087efd8bff5a01f1;
mem[686] = 144'h08c40022fda008730dac08e3f1a3fb2f0036;
mem[687] = 144'hf258f4f9077df7350eeff9460428f8c8fd33;
mem[688] = 144'hfcc3face0ec7074efbb4f05cfa740986f27c;
mem[689] = 144'h0d96f1acf45a0d16f25ff9370594f1abf660;
mem[690] = 144'hfc4cf251f1e90b2f0ad9fe98fcd4fdcf0698;
mem[691] = 144'hf76b0504f05cf748085a04ccfa48f20c003a;
mem[692] = 144'hf375f04bfd5f08780c050414fe4f09bd0ee5;
mem[693] = 144'hf346f0960e5e0758f753fef0f0a50a4ff5c7;
mem[694] = 144'hf53efa8ef343ff7af982019905a40956fb19;
mem[695] = 144'h05e500c10031fb5403bcfc5afe7b0c33f0e2;
mem[696] = 144'hfcecf071f9fefeab0bf5f3c70f860b32fd15;
mem[697] = 144'h0c69fe280d0cf1e807c40b3ffc200aacf50f;
mem[698] = 144'h04f8fc0c0ee803920d64fdc4fd16f335ffe3;
mem[699] = 144'hf7ff0df3fb3cfc7ef1d1040f0d2501bc0dc7;
mem[700] = 144'h0d7000e9f596fb3502f902c704150e26efd7;
mem[701] = 144'h0dd608a20fac0a99fc270271f0470aecfcf8;
mem[702] = 144'h02f2f4dff562f16d07cbff6dfbc60929f021;
mem[703] = 144'h0dbc02f8085ffbc6f50c06050c480ac30f39;
mem[704] = 144'hfc5b099cf8ff0999fad809210e840f51f665;
mem[705] = 144'hf4d0f9960e93ffd1095901d1006609b805f7;
mem[706] = 144'hf3a3f9b3f6190dcbfab2fc020a5106720007;
mem[707] = 144'hf5810b0cf86cf0a803830005099bff7a0bab;
mem[708] = 144'hf36f0a9608cc041b00dff3a20964f38208e6;
mem[709] = 144'hfdb8f58ef9bdf9c80b660733f1c4f8e7038d;
mem[710] = 144'hfdbb09be05de0689089bf2aa058b038ef276;
mem[711] = 144'hfe6808f6faff0d9bf345f51807660234ffae;
mem[712] = 144'h0278059ef7b7f8d8fc1c09de0a5402c4ffa7;
mem[713] = 144'h0c16f054f997f166f6a4070003bcf2e4f281;
mem[714] = 144'h04abf952fd240a93067702c8011d0be70d65;
mem[715] = 144'hff840f8af48df1d8091901650c7cf2a30c9e;
mem[716] = 144'h0a5907fefd78fec5f9b7042007420923029f;
mem[717] = 144'h08ef0722feebfcbcfea4f6a2facff591f874;
mem[718] = 144'hfb64fa3703c307e7ff0c0e1cf5ddf262f75d;
mem[719] = 144'h0885f0efffa8fe8b055b08c7f9e9f198fad0;
mem[720] = 144'h0efdf8e300c9ff130b3df864013cfd450078;
mem[721] = 144'hf44bfd290a400ec3fc6f028e03530908f97b;
mem[722] = 144'h0f4bf71f0f3401e5fdb8f2dbf49e00e70c89;
mem[723] = 144'hf79ef2a2f488f99c0dcbf508f497f52cf47c;
mem[724] = 144'hf904fab8064f09d7f2eb077cf9140970f2c3;
mem[725] = 144'hfc90f7d9081dff1a0dfcf33b05db0a81068e;
mem[726] = 144'hf73300ca052bf61cf033f261f96408c00317;
mem[727] = 144'hf97ef7e1f022fd0efbacfc45019af7fd07bb;
mem[728] = 144'h0fa00788f77f09bdf3230769f6a405b101cb;
mem[729] = 144'h087d089aff080007061df1cf0cd8f5dc09ff;
mem[730] = 144'hfb6af4a5f763f33af514f25709ea0ba90d93;
mem[731] = 144'hf2180d14fdc8f802fa4affe402b002db0d2c;
mem[732] = 144'h0a70f3d2f8510f98f861f9f509540344f52c;
mem[733] = 144'h094904c50fa7f09606380fe7f5b6f83b0874;
mem[734] = 144'hfe8bfd52f588f185f77b022a0886f7aaf0de;
mem[735] = 144'hf553ffc8f06e08fe051cfdd8fcfb025dfb8a;
mem[736] = 144'hfec804b7f7b3095c066f0f64f488005e069d;
mem[737] = 144'h026dfc460dbffdd0f4b10056fa140893fd17;
mem[738] = 144'h0078060a023efcc3095af824076704b008ce;
mem[739] = 144'hf8f2fd83f101f9890901f9bbf262fd7f0502;
mem[740] = 144'h0b9bf89b0fb0f0b0ff790c7b0fbd0bc6f5b9;
mem[741] = 144'hf7d80faef8dc0512f9f40f1ff82d00c1f0d3;
mem[742] = 144'h0e19f3060cfa01e4f7e90e0df46c01a3fc5a;
mem[743] = 144'h08000d1af90bf07ff2fbf7b601f0fdd10882;
mem[744] = 144'hf05bf790fb61fd8f07a70dae0bcd00ed0101;
mem[745] = 144'hf57801870b00f7c20478076308c2f1d4f5c3;
mem[746] = 144'h060cf3f9f5100017fa11f0f0ff88f1ccfda7;
mem[747] = 144'hf45a001e0465002dfeedfd2e0594fbf70b4e;
mem[748] = 144'h083ffaf0fa57fd700c29f43dfe8f0b68f377;
mem[749] = 144'hfc790ca20e04fd2bf7b1fa2ffad3f02df676;
mem[750] = 144'h037b0a710789f610fdc5f107f066f954f7d2;
mem[751] = 144'hf55df1b30a1af0f5f840031af3c4fe18f207;
mem[752] = 144'hf72bffc8f8dbf312052708e9fafe051f07ee;
mem[753] = 144'h07550bf80194fa060b9b05a3f901f8d2f6b0;
mem[754] = 144'h003f066802a9fe21f487fabff4cb08e5ffd5;
mem[755] = 144'hf14cf153f9420a6e0828f35cfe400b9e02f9;
mem[756] = 144'hf383f37702f9f060fa4cfe2c0f8df31df616;
mem[757] = 144'h048904f10cdc05e00f0ffd4af0abf03c00aa;
mem[758] = 144'hfc14fe8bffac03c4054900420ed3f965ff13;
mem[759] = 144'h0f7b02830b0cf2d00a0c09f00c69fcd2f9ce;
mem[760] = 144'h03e20c36f5e5f23af577f31ff43bf2f40003;
mem[761] = 144'hfeb1f09bf5d4fb99f6660637028e02010b21;
mem[762] = 144'h00aaf227f4610a15061af969fcbb08cefd1b;
mem[763] = 144'h0af3faf0f00ef2bf06340fe60ab5f1c40f50;
mem[764] = 144'h064d07b6f357069b00a40436f8ae0fb9f3c9;
mem[765] = 144'hf733f42bf46102560abd03d705fa04ba03ab;
mem[766] = 144'hfe070a810f6e0d5c036606e209ae0fa703ef;
mem[767] = 144'hfe4bf6390ee30a9e010505a6f213ff0c0bea;
mem[768] = 144'hfa86f20c03b5fd5700c605b0fb2b0b6f0c4b;
mem[769] = 144'h01690e61fefef315f3e2ff3c09cb0313f903;
mem[770] = 144'hfa660b420e6606740375fc000ad403c6085e;
mem[771] = 144'h01a503440c9af45dfa700bdcfee50501006d;
mem[772] = 144'h025ef5d0f500fcc20160fd0f0128f21bf32c;
mem[773] = 144'h04b1f3c30575fdfe0c6c096f02ef0839f84a;
mem[774] = 144'hfb7f0ec7fed3f4ddf6460f77024102e60f93;
mem[775] = 144'hfe710ae6fa1206960ff8fa24f6efffd0f64d;
mem[776] = 144'hf47f02ff020ef4a90885086efc62fc83f175;
mem[777] = 144'h03ecfae9fc220b8801480ced05f20c12f788;
mem[778] = 144'hf81009aef415fc2afe760838fb03f33a0fde;
mem[779] = 144'h0b7d0abe00400a47f5c609010826fd23ff1e;
mem[780] = 144'h09930220f2cef75803450989f74ff400090c;
mem[781] = 144'hf466fc5afa4ef612fcd2077cfad805b30e1b;
mem[782] = 144'hf0bcf628f069f097fda0061e0db5fe940b5d;
mem[783] = 144'hfbcb02a4f650084407e10c590747f442034b;
mem[784] = 144'h042c01890336f2b00b150d1b053cf135001e;
mem[785] = 144'h05deff66f30409870d800b74fd4cf38e0abb;
mem[786] = 144'hf65001e2f333f8520dc7f4ae0173000f0558;
mem[787] = 144'h0e280768f5380a1100b405b907920eccf7d3;
mem[788] = 144'h0d80fc48f42ff6b50e9dfd3e0c9ef1ed0d1d;
mem[789] = 144'h03e40a5cf954f0c00a4efdc6f13d0b380043;
mem[790] = 144'h0fb4fe4f053a0e7b0fcb0703f68ef53df53d;
mem[791] = 144'hf6c4f0230e1f0cc7046e01f30394fd0b000b;
mem[792] = 144'h09ad02d40afc00c505c3fc3af454fe4f0af1;
mem[793] = 144'hff0b03c2f2320d95fed10d700fb9f9c1f81e;
mem[794] = 144'hfb3efe960354f454f0ca08920cc108ac0ece;
mem[795] = 144'h0f99f2a8fc51fec7f35c06ad027c00410e0a;
mem[796] = 144'h0cbff6f6f55af28d0371ff390c3dfa79096e;
mem[797] = 144'hf9c306be08ba081d027d045ff5abfa39fd22;
mem[798] = 144'h0180f0e5066d07f3f8280c3e0aac04a401b2;
mem[799] = 144'hfa60fa50057ff5780baffb97059af782022c;
mem[800] = 144'h042b09abf3fc08a7f48cf8effba2f3a1fd41;
mem[801] = 144'hf34fff3bffca0b0e015efa3608ee05d80a6e;
mem[802] = 144'h0b6102070be5f0e90452fa160e88ff4f0f29;
mem[803] = 144'h092105bd0f9b0b8e04860a430646fca60f26;
mem[804] = 144'h0f4e0ac9f57202cafbad0bfbf789fe8ff189;
mem[805] = 144'hf0bc072dfa39fd24049909d6f31cf7100f23;
mem[806] = 144'hfa4af5090de2f68508050697f84afbe10e14;
mem[807] = 144'h04d7049605350a8df9acf923f6c50b58f0ed;
mem[808] = 144'hf260fd0cfe47f926f6f4ff7c0edcf1b009c4;
mem[809] = 144'hff8ef4600bbb0e2e038ff9e6f49f04a60ada;
mem[810] = 144'hf58803010eb70737fac1f2a3f87108d50a32;
mem[811] = 144'hfaecf2c6fe1b04b306d6f9a0fc92f3540fcb;
mem[812] = 144'h00660233f16cf07c0b46fcc404a008a5f17c;
mem[813] = 144'h0837fc32eff3fd1ff4c204af01d70d7af0a6;
mem[814] = 144'h097df11ef2150f3d0055f606f2c80e91fe31;
mem[815] = 144'h0b9bf084f640fd1a0acbf903ff15f4def8cc;
mem[816] = 144'hf4cb0eb705f0f848fdd3086e0fb506390728;
mem[817] = 144'h0084fe9bf4f7038ff0aafe96fd8e068efddf;
mem[818] = 144'hf89200fd0c860e55f187f8fff26af386f3bf;
mem[819] = 144'hf7b9f1f3f43301b1005c0e46010ffd2e0d51;
mem[820] = 144'h0cf0085ff21c0a53f0d800deff4f0c240d1e;
mem[821] = 144'hf7f606dc06ef0ae40ab8ff82fb8efe640a2e;
mem[822] = 144'h0c8d02a9fa750c0bfa82f967f2e70cddfec9;
mem[823] = 144'hf526f84ef054ff850b5409cb08790d14fdb9;
mem[824] = 144'hfa8ef2810081fe68011e01f9f27506f1f1af;
mem[825] = 144'h0603f075f304f05ef610feedfa5bf726f7da;
mem[826] = 144'h05fdfaabf5aaf3280911f9c5069df1100513;
mem[827] = 144'hfbcc03e5f406f67af4f1f911f15df51af55b;
mem[828] = 144'hf775fbaf0c220fd80030f69cf0d00295f15a;
mem[829] = 144'hf1ba06cc0e04ff99fd7e02dc0881fd1f0021;
mem[830] = 144'h01cbfa34fdd5f29e0b4c0cf7081a0523f826;
mem[831] = 144'h0144f7060db10d50018ffbd00f68fce5086a;
mem[832] = 144'hf053f8c4003703fdf448f290fbf008170913;
mem[833] = 144'h04780994ff7af2cff250f9e509bb0c57f3f4;
mem[834] = 144'h013c0b66f6d50fe006580a3e0de00d510bd0;
mem[835] = 144'h064305a5fef4f094052e042df69a08ef04dd;
mem[836] = 144'hf19f0f97fc0207f807aaf4160d0afb21f3e7;
mem[837] = 144'h06c601b1f5d70d52f182013ff03f0c650b7a;
mem[838] = 144'hfbd40e8af0bef76d01510e3d05b6fd220e26;
mem[839] = 144'h0667072a078cf8b50ddcf5e30750059502a0;
mem[840] = 144'hf81b0725070e0956038ef3a408abf9890c8e;
mem[841] = 144'hf109026400930da608c4f45af3bbf10ff6ab;
mem[842] = 144'hf5f3f6c4f1d00847fd34f68cfec3fce5f07a;
mem[843] = 144'hf9f0f43df7ee0c17007c0263f18e0ad50d5d;
mem[844] = 144'hf0020bebfa79fe850731f71bfc3901cef5c3;
mem[845] = 144'hf3edf47bfeb103d80222fa5e0121f84ff0b4;
mem[846] = 144'hfcc0fc080ba50adf0c37f22aff2b05f50f9e;
mem[847] = 144'hf25e02bc0d6405a70e36000ef8750b240373;
mem[848] = 144'hf860f39efb0df4a4f36bfa4bfb84f6b6f9e9;
mem[849] = 144'hf549fb970c9cf898f3f503c4f315ff720ea7;
mem[850] = 144'h0182fe22f54408f1f839fae7fb74fdbe020f;
mem[851] = 144'hf06cf9d2fbd1003af7630062f4f20cdbf389;
mem[852] = 144'hfd3206c0073e0dbbfa65f6c4053dfdf9fb51;
mem[853] = 144'h0751fbfafde8028f02ecf058fed1f2e20caf;
mem[854] = 144'hefe30b0908bdfea4ff43fcf60e070a83fa93;
mem[855] = 144'h0243faa6fc2bfed1f200f08d057efc14f231;
mem[856] = 144'hf2290b2506fd0a640b86f2d408980fb90800;
mem[857] = 144'hf2b203a600a9f8c9f9e1f2dff2d3046808a8;
mem[858] = 144'h0ba201c90641067a07bcf0520351f619fc41;
mem[859] = 144'h0fcb0f55ffd50a9400b9f455f99b0901fc2b;
mem[860] = 144'hfbf1f3c404e704d20d03f7a30bf407feff22;
mem[861] = 144'hf7020e92fed209be0004f177f1be0294f822;
mem[862] = 144'h0699099d0dd40ed005a5f264f922feb6ffa5;
mem[863] = 144'hffd40199f980f10e0feb03870373f21d00a3;
mem[864] = 144'h003a031e083bf80dfce9012405f6fd6c0c42;
mem[865] = 144'h04f00783f09cf6d304e40884fbd30c4c0ef6;
mem[866] = 144'h0ed3fc4404ad0fa9061b0be7f224fda9f3d8;
mem[867] = 144'h0897fb25050a06d60f7101cafcdf056b0077;
mem[868] = 144'hf9f9fb08fc7300c9054af562fdf1f432f76a;
mem[869] = 144'h0c8bfb1efbaa0aee0fc1035ef3bcffe1f994;
mem[870] = 144'h0859f2c2f2b70cf3f6eff32ef4e70f260c72;
mem[871] = 144'hf919f4c40ff7067f0759fc31feee0be405d3;
mem[872] = 144'hf8b7fafff1c70279f0e30186fa15f2b40d55;
mem[873] = 144'hf01303300132f302f26e014302870143f9a0;
mem[874] = 144'hfb5c0c03f3ab0c17fdad04b70d350317fca7;
mem[875] = 144'hf519f28df89bf35ffd3f082c0788fc8e0d49;
mem[876] = 144'h019ef28b019c090b0cc7085efc57f979ff7a;
mem[877] = 144'hf1040eadfd3cf4f60b250bf80e6ef5d8f55a;
mem[878] = 144'h057d0e9e09c9f7200543fd5afdb3045807b2;
mem[879] = 144'hfa2108df0086f22f06b506ecf79cfec5f300;
mem[880] = 144'h08210047f6160270fbda0deffc63fcfc0ab5;
mem[881] = 144'hf6150e0cf4fefa1402fc09edf8c6070cf8bb;
mem[882] = 144'hf87302e0f590ff8bfb8df85f0eb7f0db0ed7;
mem[883] = 144'hfa7f072b0bf0062ef2a10f93fdeff56fff64;
mem[884] = 144'hfd8b0133f1270126ffebfb590b5304e801f1;
mem[885] = 144'h010ef289f69bfb61f811f72c06d5f73e0c25;
mem[886] = 144'hfd830b400123029d0932f140055501d3f0fa;
mem[887] = 144'hf0dffb52f64508440980f3e8f7f6f57a0bb5;
mem[888] = 144'h001d0bbdfca508f001e7f2d9fcf2f048f13c;
mem[889] = 144'h0a1cfa84ffbf09f80357f42efee60fa808c5;
mem[890] = 144'h070ffe83f83b0aeb05b3066404b304cff2a6;
mem[891] = 144'h0f6c0232ff22f54ef3d1f02df99a0a0ef0f1;
mem[892] = 144'hfdde0e2b0ce9ff5e0cc30bb80b30f9150914;
mem[893] = 144'hfe140426f0370fba087c056ef1b20a420a55;
mem[894] = 144'h04b408e6085cf1e40e8c064bfd89f1dc007c;
mem[895] = 144'hf68b0ca3f436015400eef08001dbf0f8f8a6;
mem[896] = 144'hf9f90e4209def03ffb13ff45f5a6f5b3fd14;
mem[897] = 144'hf2220a8c07fdf906f8fc07460ab6f6ea0568;
mem[898] = 144'hf847f993f3acf408014308ae0497002d0abd;
mem[899] = 144'hfa46f364f9630c7dfd1203f80f22fa32f22c;
mem[900] = 144'h0d4607d0f02e05480b6cfbaafcac01330258;
mem[901] = 144'hf5e5f69000dc0b36f34d05f60542f371f823;
mem[902] = 144'hf41f0e1f098bf1220446fc9508ff05dc06c8;
mem[903] = 144'hf79af047f4c00f94f249f095f65ff332f178;
mem[904] = 144'hfc820a2e0c76fb4cf2c2f482017af6370054;
mem[905] = 144'h036609f8019c0437f80bfa920c5ffd330c71;
mem[906] = 144'h0ac80a52f04dfa560cc108bf04c7ffd80fd0;
mem[907] = 144'hf3a60486f6aaf6fb013ef07bfb2009d607ef;
mem[908] = 144'h032802e1fd460a8a066ff59d0add0bf3fbf1;
mem[909] = 144'h0135fa90f696fc4e0d070e27ff31057afd70;
mem[910] = 144'hf25c032dfa89003afea3f2b9ff1a0c39f22a;
mem[911] = 144'h05c7ff61f36503ba08e7feedf986f2e2f27e;
mem[912] = 144'hfd1b0e270e6cf16d075af5ec0d1efda608c2;
mem[913] = 144'h09620d48021afe0ff3870c5c03490477f88b;
mem[914] = 144'hf9abf334fb73fea4f6e5033ffd360ea0f1d3;
mem[915] = 144'h0844f7f9f8b106330f490b290d8cf8aafc6f;
mem[916] = 144'hf91b0db504f50ba607b801a5fefe074df9a0;
mem[917] = 144'h083ff28a0a880c68f78a004901bffe5df624;
mem[918] = 144'h0b340f80014df8a4083a03040cd5014e0b2c;
mem[919] = 144'h04d8effd097e06cdfea0fd1701a1f46df23c;
mem[920] = 144'hf008f5e80199f0d8fabc0c57fda809a7030a;
mem[921] = 144'hfdb0fc45f5f7020b0673fac6f4ab0e2ff5ef;
mem[922] = 144'h0b5a0354f286f30108930ac70e41f80bfcc0;
mem[923] = 144'hf6a7ff39042d0f32f2e6fabc018d0722f58f;
mem[924] = 144'hf2adfce2fdacfac10ec70bccfd0d0e20fafa;
mem[925] = 144'hf789f8f5027201270010f3b60828fc26f61b;
mem[926] = 144'hf4e709450df80ee00a02f35f02bbfc9ef81d;
mem[927] = 144'h04c90e9f0219fca0f030f0b3f3faf39af116;
mem[928] = 144'hf7ccf144f58c0d81f99304360b6803b2fcfd;
mem[929] = 144'hf9ac09a201dc0e4cff42efde0e3ef8670144;
mem[930] = 144'h01cefbc9fcd307a70cc7f0710310f8a9f8b1;
mem[931] = 144'hfc17fe05f25f0dcbff7cffa9f9a8f75e09be;
mem[932] = 144'h0265f41b0815f5a6fcb1f431fe5bf43a08be;
mem[933] = 144'h03b5081fff0403f4fa1df614020ff0d5f5d4;
mem[934] = 144'hfed809d609a9f7e8079df055004007dcf93d;
mem[935] = 144'hf7ebfc3d0ee0fe6405ce0b3408a2fa47fbca;
mem[936] = 144'hf3fc04effcc00b300851f846f3acfed9f11f;
mem[937] = 144'h0de80c19fd2cefcb0dd1fff5f2660f910aaa;
mem[938] = 144'h0e830671fc3e05f5fe9305730fb0f72bfda2;
mem[939] = 144'h04fa0b29047e07500e550b54f603011ff5ed;
mem[940] = 144'hfdd10f9b0805ff8b05a0fa27ff94004306d6;
mem[941] = 144'hff0504f101ca023fffbcf506f6c2fe3609c4;
mem[942] = 144'h018cff87f5eefab5ffed0add02270ee20369;
mem[943] = 144'hf01a07b7043cfedcf2a9f842fb92fa73f719;
mem[944] = 144'h07a4fc5ef4a00686f9db00a30dcf0de9f56f;
mem[945] = 144'hf5c3fe170be8fc230ce4fb61049b055af47b;
mem[946] = 144'hfc08f6dff2a40583fbc40636fae8078efce6;
mem[947] = 144'hf6d402a5f5ecf0260370f0670b7906640929;
mem[948] = 144'h09cff712f21f063e00530681fa590c99f065;
mem[949] = 144'h0dbff1f90402fcba01a70aa4feb3f73f0b7e;
mem[950] = 144'hf02ef7c8f9f3f6a4f3d6f974fc0c046c03a6;
mem[951] = 144'hfeac0c230d410036f276f57501f309e1f5b5;
mem[952] = 144'h0d20f27f0f57fab501960b0d083bf9c5f2ed;
mem[953] = 144'hf097efe6f662f95506f40559fa4ef6230b9d;
mem[954] = 144'h0bc3f3b10c17f27cfdd005b6049ef7be0cd2;
mem[955] = 144'hf897fc220fb1f88e0c81fd050294f09df46d;
mem[956] = 144'h0eba0adbfdc4f73d0071f3480d3af484f538;
mem[957] = 144'h01390d8bfc45fcc2fb6bfb68fdadf0c303e6;
mem[958] = 144'h098d004ff16dfa7a0ee5fc41fac40487f087;
mem[959] = 144'h0c170526f4f2fe8b060904780297f7620ed8;
mem[960] = 144'hfa780da6fb4bfd28f140ff6703a7055eff40;
mem[961] = 144'h0cbafa7c0ad4f1bdf27f0d85f33e0e370604;
mem[962] = 144'hf7c3048b05cd0bf5f284f076f6ecf3b303ff;
mem[963] = 144'h01fff9cc084e0a36f050f7c001e1f9e2f3d4;
mem[964] = 144'h06fffa7ffadbf60802aefb5c0bddfea7f88c;
mem[965] = 144'hff8f0290f62cf808f977f315fbd3ffb2fe38;
mem[966] = 144'h0e03f87dfcb0059e05d8fb11080df4a90f5e;
mem[967] = 144'h09e40e0c0881fb580e22f37e00170501f1f7;
mem[968] = 144'hf8ad047408d7fca8f4a6f1200515f90f0f0d;
mem[969] = 144'hf5ba0a0af5a00c200145f06ff67e0baf0767;
mem[970] = 144'hfcc7f9700dc0004ef01509fc067bfd960ef9;
mem[971] = 144'hfa3ef1ecf893fc82f705076ff148fd86094b;
mem[972] = 144'hf77f04f405fafa8e088ff8b40ce7f04cf584;
mem[973] = 144'h07fdfaec0c0df88405800f9d0d8bfe43f766;
mem[974] = 144'hf1f7f9100deef969ff9bf8acfd4dfb190cb4;
mem[975] = 144'hf57b0a07f1610d3d099700e003050a80f957;
mem[976] = 144'h058c0fd5030e09aef615fa68f832f5360788;
mem[977] = 144'hf4b9f3c1062b0d21f27b0027040b02ed0e3a;
mem[978] = 144'h058908d801800829f0fd05cbf135089e0d69;
mem[979] = 144'hf70ffdef0d1bf1160897019a01690f29fd2e;
mem[980] = 144'h0cd6fad2ffeaf65c004304b40c43f3380dd3;
mem[981] = 144'hfb56f90c0feb0fd30699f8abf11ffb03fc5f;
mem[982] = 144'hfc13f35eff0701af07e90605fe7e0acd003c;
mem[983] = 144'hf9effa96fddbff80f3d9f4490deef796fa73;
mem[984] = 144'h080f01ff0e6f08b10c41010d0b800f5efa17;
mem[985] = 144'hfd9efb0e0548fe070cbf07acf6c60657fd4b;
mem[986] = 144'hf75905d6f5f2fdf80b68f01cf6fef98f0750;
mem[987] = 144'hfcd5f5f9f1c20374f2bdf719099f091df35d;
mem[988] = 144'h052c0a88f850fb9808f1f978fd6df465f873;
mem[989] = 144'h0702fd7d0252040af918f625f1550b3ef08a;
mem[990] = 144'hfa86fe70013a0d1f06eaff840ee8f98701f2;
mem[991] = 144'h0e96faff0ce6f554033ef445f76209c3fece;
mem[992] = 144'hf7c00969fd44098109fef582f0b4f738fc27;
mem[993] = 144'h077ffe45f9cb0151f292f8080298f98b04cb;
mem[994] = 144'hf81efd860f8903b303fa0c03f4aa084cfd43;
mem[995] = 144'hf529f9cf049000780798f3060ae50b8a0985;
mem[996] = 144'hf1c50bb9f9e808990757fd60faf9fcca0ac1;
mem[997] = 144'h09c10090f0070457fdeafe370b7a02c40a98;
mem[998] = 144'h0badf942f839f64cfb56fa8a0209f3f409c1;
mem[999] = 144'hf58cfc40f1b006a6066ff499fdad067d0b82;
mem[1000] = 144'h0f040d1903610e28f21b07030dae08340276;
mem[1001] = 144'hf6daf9bd0353f732079f06ddf106f720ff04;
mem[1002] = 144'hfed00802000bf8e7fdb80bf3f5e0f2680051;
mem[1003] = 144'h01d9fc11f8c102c805e50590fb77001d092d;
mem[1004] = 144'hf4baf8cef27c00b5fad906ca058dfb550f65;
mem[1005] = 144'h03ff013e0dcb06acfbb3fd27fc5ff9dffac5;
mem[1006] = 144'h07560be20e78f2f5f2880836091a0c660d42;
mem[1007] = 144'hf229fce5f77207af01960a7c0d010f9805c2;
mem[1008] = 144'h0614fbb001300b370f50f019fbe50546f510;
mem[1009] = 144'h0e09f7c3f32cf8d2fe5ef4d2f405fbbff5fd;
mem[1010] = 144'h0ea603ccf699f8cb0dccfd9bfbda012406a4;
mem[1011] = 144'hfcb70d4d008e04bef6d7ff14092b03d5f816;
mem[1012] = 144'h0b85059f058100f10750083c0e860bc8f0bb;
mem[1013] = 144'hfa0d0ef2037b08240aea02250e8af761f69b;
mem[1014] = 144'h0bb6f51f08df0f60f5ecf40efa5905f8060d;
mem[1015] = 144'h01b6ff620e8309fa09a1008c07ff084c0309;
mem[1016] = 144'h022d0a49f7b0f3ddfa63effdfed6f401f52e;
mem[1017] = 144'h0604f93ef0e00734ff58f7ad0f3a02fa0477;
mem[1018] = 144'hfe33013df41f0625068efe18f8e3f637002e;
mem[1019] = 144'hf36907bf0dd2f7bb046b0d12f79f0379f6eb;
mem[1020] = 144'hf9ddf3adf8f60e40f3b8f310f50ef3faf2a9;
mem[1021] = 144'hfe0605c002d2f9e8ff8e088ff8510cd6fba0;
mem[1022] = 144'h06ebf789fc67f996fdacfbcd0fd6029af0b1;
mem[1023] = 144'h043cfb0fff07023107ae0a1e04bb0365f65f;
mem[1024] = 144'hf75402bbffd907f4fc2505f106e80bfffe56;
mem[1025] = 144'h03d8f3b809eb00b20147f5ed06ec0e77fa66;
mem[1026] = 144'hffedf8c60d5cfab0fa3304110c0ef5490edb;
mem[1027] = 144'hf0a504fa066e0806fcb5f59301200c1e02cc;
mem[1028] = 144'hf03ff08b09def015f636f7c6f9e90ea30ee6;
mem[1029] = 144'h0f3f05b60a2a0c12f7c6f33e0ce70c450cb8;
mem[1030] = 144'hf07b0770ffcff0e70254010ef8960e16f12c;
mem[1031] = 144'hf70503a8f4c5077b0090fffcfd2d00fefd3a;
mem[1032] = 144'hff46fb5b02150508f0ad08ff0a3c03df06d8;
mem[1033] = 144'hf9daf7f10f44f51d025e0e50f6cef06a07f5;
mem[1034] = 144'hff5a06fdfaa50224fb650a300479f5700b4c;
mem[1035] = 144'hf424f6b40176f961014a09aa01cefea3fbd8;
mem[1036] = 144'hf20ff9e90e88f5af01edfa7cefe00ccc0b62;
mem[1037] = 144'h0194f938011ff4550406fdba08d7fc1b09a2;
mem[1038] = 144'hf757fff1097ffc52071d01bcf0c2f4eb0854;
mem[1039] = 144'h027801a7fe52f9ff0c7ffe4cf1b3099e0248;
mem[1040] = 144'h0380fcacfd790ba10749fd7f07470bb003ff;
mem[1041] = 144'h01b6086df25d0ee5f550f60aff4301aafaf3;
mem[1042] = 144'hfd73ff47053a0ab507cf02b0fe010dbefde8;
mem[1043] = 144'hfd6af5a6f15ff8d8f83dfa64effaf9d0f128;
mem[1044] = 144'h06f8008a05a70e77fe63f6050dccf0adfcb8;
mem[1045] = 144'hfc07fccefd1dfece0a43f38408280225fead;
mem[1046] = 144'h0bf3fe10040404aff8600cd6075bfe57f390;
mem[1047] = 144'hf62bf378f47c0e2301bd01e908d2f4f90002;
mem[1048] = 144'hf3c0084106e5f254f8e6fd2ef2d2fe94f0b6;
mem[1049] = 144'hfe510a29f7c101e70c80f388fcb906c60ce7;
mem[1050] = 144'hf595feba02a3fff708ef0a7803a0f299fd16;
mem[1051] = 144'hf24ffe1501800a18f860038f03f3037ef392;
mem[1052] = 144'hf7ddfb5b0b49f4f0f6f20b7d02c90f2dfc3e;
mem[1053] = 144'hf6a2fad1fa37f961ff6205490f2dfd3a00d3;
mem[1054] = 144'h01f70270f1f9fe92fafef34ff18ef05c0874;
mem[1055] = 144'hf01bf3880fa0f22ef34d0ae80ed4075af1bf;
mem[1056] = 144'hffc6000df6dafa6c0c300e62f5cc0d31076d;
mem[1057] = 144'hfa580076f959064ef1f6facafe85ff5a09dd;
mem[1058] = 144'h0229f9d707aafc57f93df7440468f673041e;
mem[1059] = 144'hf01504930c5f033ef27cf36dfbb203fe05cf;
mem[1060] = 144'h06bf00640dc80c0b0098f4e3f52e0e3d007c;
mem[1061] = 144'hf2d1f31f0c72f8bf0a66f07cf8f90a60f538;
mem[1062] = 144'h0baa07b80064f30bfc87f8fff029f3900f95;
mem[1063] = 144'hf9c4f9a006b5fb080d64fe1ffcd4f75cfaff;
mem[1064] = 144'h016407450196fda7f688f602f95f0569fad0;
mem[1065] = 144'hf479f7d3f84504c6f154f43ff1c20084f88f;
mem[1066] = 144'hfbfcf12cf692f18303590be40bb2044a023e;
mem[1067] = 144'hf594f61c07f10df2f00801def98105caeff1;
mem[1068] = 144'hfdc3f578f0b100dafb0200b00961f662f867;
mem[1069] = 144'hf214f8740fb0fbeb00340f430c3c0537f5ad;
mem[1070] = 144'h09f5f97ff9a3f36f06bc0f6bff940eb5f926;
mem[1071] = 144'hfea90a62f7520c4bf28ff2d70e9808970500;
mem[1072] = 144'hf924f945fbeafcadf06c0b29f2f404fdf623;
mem[1073] = 144'hfd43f77209c30e3bf74cf981fdcf09c50ad7;
mem[1074] = 144'h039b0a75fc1cf292f3fa091bfc66f0a10cd9;
mem[1075] = 144'hf16ff12105860c70f70bfdb4fdf404490a75;
mem[1076] = 144'hf59efcac04720be9f4c50fb80e7e0d800769;
mem[1077] = 144'hf0a2fd430060ff2bf829fd9cfa8df55ff899;
mem[1078] = 144'hf36e0ff90b06fc3ffa4400e204bef1f8f84e;
mem[1079] = 144'h04ce09690e42055f0ed4fd5ffb39f62bf41f;
mem[1080] = 144'h065ff28efc720e2708ac0567f28806a1ff81;
mem[1081] = 144'h09e2fce9093af14ff414f4c3fe460761fbaf;
mem[1082] = 144'hfbb9f19cfba10d350157f8c9f8f1f743f816;
mem[1083] = 144'hf5f2f9440326f2660292fbecff1df7ed0d62;
mem[1084] = 144'h06540e29fe580e8df05efbd10afaf2860925;
mem[1085] = 144'hf40708c80c2e068606caf37bf373f931048e;
mem[1086] = 144'hf3abf43f0630045aff63080d09310072003c;
mem[1087] = 144'h065cf568f46908c3074cfdd10aff00ddf1a7;
mem[1088] = 144'hf7cbf5710b4bf7d3074af347f560f561fbf9;
mem[1089] = 144'hff04ff70fb3bf7c3f2dd0daff1e90acb0c69;
mem[1090] = {16'h04a9, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1091] = {16'h0218, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1092] = {16'h01e8, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1093] = {16'h08fe, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1094] = {16'hf397, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1095] = {16'hf5b6, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1096] = {16'hf8bf, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1097] = {16'h0707, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1098] = {16'h0b8f, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1099] = {16'h015b, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule