`timescale 1ns/1ns

module wt_mem7 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h0f8205bff4741c19ec0b1a241f2feb2af27c;
mem[1] = 144'heb0505c40a1019a1ebc5f8ef060018bd03a9;
mem[2] = 144'h032aed48eec007d5f345160f0591fe28ec7f;
mem[3] = 144'heca800000708e1f4feb407900f9d19e616fa;
mem[4] = 144'h0c6f0c27e7e409e20a691fa301c0eb48ea95;
mem[5] = 144'hf0a6fbe917cae9b201a300ddf1d3fd211c2c;
mem[6] = 144'hf986ef7a0263150b06bc178714c804cbf08d;
mem[7] = 144'h0ffb12900af6f7ed1cacfc0ced9bf4a0150e;
mem[8] = 144'hed3de1f4e2ff030d0740ff3e07ecf71cec50;
mem[9] = 144'h0286f26210d90d26fa85145b1fe3fdbbe662;
mem[10] = 144'he3f106e7e82f11ee0f71032cf59be6b5ff0e;
mem[11] = 144'hff35f178fb7e1137e262fce9f9580b170711;
mem[12] = 144'h0f82e7fbf44dfb25e18d09d5fb78f28f1d6b;
mem[13] = 144'h17791fcf06b30865ee5af8cdf6ba09cae91e;
mem[14] = 144'h0ad8f53ef2d41e890a660bb7105befae01d0;
mem[15] = 144'h13e5e9051acefefaf9090dac19131b36076e;
mem[16] = 144'he1a20a95e842e64fef1cf0cd1f76f975efeb;
mem[17] = 144'h016614c80581f80815f2177f1bb9f7761bb8;
mem[18] = 144'hf9291ba81498004e0d1ee8b70981f915e443;
mem[19] = 144'hf89ce304e1720599eeca17d8fd651591e50e;
mem[20] = 144'hfb95fb1c0d44f065e75cefb9f2a6ff351241;
mem[21] = 144'h1bdeeb3ce04b1412f6daf4400e39ebe90cad;
mem[22] = 144'h04f709231dfbe405ede515d8ff971541ffed;
mem[23] = 144'hfe61e1e8fcbf19e6e331f836033013481226;
mem[24] = 144'he134fe0e09a11341ef5eea1ae8dcf692f1bc;
mem[25] = 144'hea01fb18eb6c0d58181408c80488f90c0868;
mem[26] = 144'hf863e94ef353f7a9eb95107e06b5e634ee8b;
mem[27] = 144'h1aa7e9d6ff68e34515a41f9b05e5ea98f665;
mem[28] = 144'he8edfc1cf34907431585fe9ff081ebf4f506;
mem[29] = 144'h0813066de22aeea2063f00b504dffc49f9b9;
mem[30] = 144'hf3bf1293f4afea3ff1cb155216eeef3614f3;
mem[31] = 144'he8caef2916e61281ef990c82e61de6c90eea;
mem[32] = 144'hea4c03a01aeae09c18b5e99cf29ae386164b;
mem[33] = 144'h183de2aaee51e5a810ba0c04fdc10d0003db;
mem[34] = 144'h13e9e581fb2fdffaf0aaf5fee014e15b02a8;
mem[35] = 144'he61a0574fbc5f68c0abde8f505d509541009;
mem[36] = 144'heb34f11d0d53ec37032c0afa06ec1b531cc0;
mem[37] = 144'hfa4ee84af118ff9a17271750e7900629e39e;
mem[38] = 144'hff421b03eef2fe7af85c0b50ff8ee759156f;
mem[39] = 144'he7d2fa800a27eabcff19e0aae010ea2fe78b;
mem[40] = 144'he375f7f818be019013370d31e6e7eed3f820;
mem[41] = 144'h1929ff6ef229fd77e40bf0f8036a19670627;
mem[42] = 144'hf943ff42eba9fea8f13e16f8041e1f51e1bb;
mem[43] = 144'h13cae37800b5ebf406f8e192efd011ad1f1f;
mem[44] = 144'h082f03df0a2df660173019adf5d3ed61ed38;
mem[45] = 144'h0e1a03e11c2d0766142017e112840544009c;
mem[46] = 144'h0c791945f1d7dfecf3fee6b0f7ed0620f7d1;
mem[47] = 144'h14ace2d6f3c41bb6044aff25f9990f9cedb7;
mem[48] = 144'hf0fd14ff0cf5ed06135015f50672120410ce;
mem[49] = 144'hf73ef604ed240e171cf310e3166a1c7a0735;
mem[50] = 144'he56d19e4f36000fb0e100c4e15b9f84c185d;
mem[51] = 144'h07b401e7f722e1aff4cbe8a8f46a065f1a8b;
mem[52] = 144'h1d900dace4b8fc7d0b04f0bb06dbed5816dc;
mem[53] = 144'h051a0182e92efe65ee5209d613970d6308a8;
mem[54] = 144'h1afce84d156dff771089f0ad15721b4fedbb;
mem[55] = 144'h1addf07a1065f4751828e1e616c1ebe708e1;
mem[56] = 144'hec37ebc215b50c0de2ece785e33818a5fa3b;
mem[57] = 144'h08dc09c9f5b9f8a3f86a1acd1101f333fd33;
mem[58] = 144'hf57cfd8d0abf122be82514d0ff24185a0942;
mem[59] = 144'he690f84ff207fef4187de2d7faccfa95edbe;
mem[60] = 144'he584e80ae1021ca5e0b808c9e0e3ed8700e7;
mem[61] = 144'h1b690b64f97501ab1acff3ea07fae9ac0c69;
mem[62] = 144'he9a6e3bb0eecec51f8e9e69212c4f33012ce;
mem[63] = 144'h15f7e5f91222f2d01311080be1cd0d931508;
mem[64] = 144'h03ab17ef16440b6b1c531a5de5e2e622e0f2;
mem[65] = 144'hfa3fe8be0029f72e19c012831202f28e0ba5;
mem[66] = 144'hef72fb34ebebe0871382f7e813a20f8efe62;
mem[67] = 144'hed4aec89e347f734feeb03aaec1a1216ea8d;
mem[68] = 144'h0d7806bef4fbe9c7008dee2517a81aed04ab;
mem[69] = 144'heca0e013f7a7ec01effd07da01dd030d1d8c;
mem[70] = 144'hfc25024d0f57ff44ec0301241d6414c81344;
mem[71] = 144'hfe5de8d5ffcbee8815111ed6f7e3fe4b0fad;
mem[72] = 144'hf5bd01270104066a0a2ced290d42008c0d24;
mem[73] = 144'hf9140e81fe5ae29a09f0e0d01c3109cde24e;
mem[74] = 144'hfb0cf55b1edef53112e0eea1fb440a5e13ce;
mem[75] = 144'hf74114a8e1260a24f0021c450800180b0d68;
mem[76] = 144'he54d1266e1e2182f06ee13921a24fd4fe7ce;
mem[77] = 144'h122902b70d2314c51630eef2f5a4f1ebffd4;
mem[78] = 144'heef815be1a0f1cfc02ca19b6192ff8371e15;
mem[79] = 144'h05630c541a87ecdb112f1eaee84fe59cf662;
mem[80] = 144'h152f15150478f23cf27e0c52e754fc0ae181;
mem[81] = 144'h013502ed04851c4eea1d05a3e18a15b5f005;
mem[82] = 144'he1a70752ed5cf7dc002ee9bf185fe93ce6cd;
mem[83] = 144'he61ef31ef42dea5de9d50f8eece3e01e002a;
mem[84] = 144'h1ec7117be186122cf4dcf879ea051f791f67;
mem[85] = 144'h1c010e621033e6b505fe13a2e634eece06e7;
mem[86] = 144'hef8308d8e1661ec91104f0e5fa8a04ebffb9;
mem[87] = 144'hfe87fec21347e2c2f41feb7a14d4f05303ea;
mem[88] = 144'h03110cb3194fe34a19d11dc9ef7cf38211d8;
mem[89] = 144'hefe2f90fe829ee27f20e09cce0e119aae5a1;
mem[90] = 144'hf332ede7f3e5007f078104ebef141745e262;
mem[91] = 144'h04620f8d196a0888ebd012c6e1d105d1ee11;
mem[92] = 144'he55c13b5fc4be7f8fe86eecae43d1d59ee9b;
mem[93] = 144'hea9e0e3efe450b19f3021bbcfce612590015;
mem[94] = 144'hffbe0106e135f57d12c01244177aed4bee4f;
mem[95] = 144'he3d002e71221fbd60171fba8034a03e6034d;
mem[96] = 144'hf2ffe6d2e09ef21df478032bfd50f61701c5;
mem[97] = 144'h1507138e0607e7b5169b0c18f0cc12c80148;
mem[98] = 144'h162efc9501f61274fbc7f691ea3ee4601890;
mem[99] = 144'he4001e72f4251930f3c400eb066cf89c0209;
mem[100] = 144'h1d97f8aee0750133fd1c1a091a5e0380e37e;
mem[101] = 144'hf12707cc072c1c36ead0e21a1a8de05f0aa1;
mem[102] = 144'h13d1e290098b1c7b071a079a1ab2ff87177f;
mem[103] = 144'hf835e430fb78f31902eafc2eff0d0390e94e;
mem[104] = 144'he5421172ee180ca6ed120166ff7a0642f4c5;
mem[105] = 144'he8af04b1e0d7f297f990f9f9fc9d1ec91286;
mem[106] = 144'h1128e038eeb4e2200420fa130848ff751e62;
mem[107] = 144'hf142ff6c0e99056ffe27f5b4fe73eda9faf5;
mem[108] = 144'hf7a0ebde0c4c0f740cbe1c72f6fe19d413d5;
mem[109] = 144'h12d8084fe5c5075e1a8af235f44610c506c0;
mem[110] = 144'hef2df2540fd9000c0c781fab067505801be9;
mem[111] = 144'h14f2ef51013cea5611dbf1abe0b5fed01872;
mem[112] = 144'h12a3ee30e8dd175de1410344ec31104b0194;
mem[113] = 144'hfb17164bf3590e16e13e01c2f5c601880292;
mem[114] = 144'he0d4e0c2e581fca00d620949e5ab020ffc7d;
mem[115] = 144'he1a6ea94ff89fc30e861e7bceed40b0a07f0;
mem[116] = 144'hf9bbed0c136dfaadf300e7eeeef70488e572;
mem[117] = 144'he2a4f7a9ef2de83e0a6c185e0e4b02a11af9;
mem[118] = 144'hfc1f1bfd18d6e9c30e14fa9c024aeef5ffd1;
mem[119] = 144'h1fc817b806d0fe47e419fa7d179b1da10895;
mem[120] = 144'hf6250a8afc97119be84409fb036a005a1ccf;
mem[121] = 144'h14b3f895fa3ee27806a6fae903790272e403;
mem[122] = 144'h1547e082ff74120c1577ea6ce4fdfb4f14b3;
mem[123] = 144'hf1eb0495f1bbe2beebf5e06effb0fef9f232;
mem[124] = 144'h1c65eae4f47bf1eefb37ead3f1151b28f6c1;
mem[125] = 144'h0020edbff7430b01f2f80dade630e5ad1193;
mem[126] = 144'h0e091734e525e3d602a51bcc122bf0e8e5cc;
mem[127] = 144'h1eefe73d1c84f2b9145c01d307f0e5c3e829;
mem[128] = 144'he3deecd8004affd3fb63eed1e33a0358f9a1;
mem[129] = 144'he7b1170e0fa61b48eba1e55501bff9830c62;
mem[130] = 144'h0357e259ef5ae662038e1bbcf41f0fb30ac8;
mem[131] = 144'hf56711c4e3900af0f603f12d0446e2881dbc;
mem[132] = 144'hebf6f8bfef86e6f30bb7e2e20be8eedb1d85;
mem[133] = 144'h0962f3071b60f5680ed91f08fd431858fcb8;
mem[134] = 144'h18e2114319961faa060bf463efece9d71d8e;
mem[135] = 144'h0a4bea6a0880f617f1871de00725ea8a082c;
mem[136] = 144'h1baef2deff2d14620818ecb9fc4beadee18c;
mem[137] = 144'he8cef792ed9f090ee633ed44f4b0e2c2f128;
mem[138] = 144'h148201270d2d0d5ffd49f7b517ef12c9f34c;
mem[139] = 144'hfc0ef7a60c28040b1cd9ed81f5000d611bad;
mem[140] = 144'hebb0efb9e70ef80aed3cec621a0e0aca17d4;
mem[141] = 144'h0b7b00d80820f49e10980be01046e99c1912;
mem[142] = 144'hfc9aeddceb71e499fdbf03770bf8eb38f52e;
mem[143] = 144'he7d5130be3bcfa8cf31dea2ae6af1957f674;
mem[144] = 144'h09de15ef0f74f961f99c03c4e73d15dde095;
mem[145] = 144'h0fb2f0aeea01fce004691678f1dfe07efb76;
mem[146] = 144'he7a9f985089d1393f052e5f906df157d0e9b;
mem[147] = 144'h03a3f5d9e614ed780a701b310340fbd3046d;
mem[148] = 144'hf8ebe42912b908691b2f0c2208f41316f9f3;
mem[149] = 144'hf8bfe388f8711383e916098ef156f8380888;
mem[150] = 144'he6aef931f2d208210e42f33c120b0df6e4a9;
mem[151] = 144'he3d7f9ad01a5150bf6c5e6e216250472164a;
mem[152] = 144'h16251db513d218d5e18be5e30ac613d0f524;
mem[153] = 144'he6a20e831263f6bbf7d112c917c31b28f0e8;
mem[154] = 144'hf189f66ffb2f11caeb7f068bf1f7f90104d1;
mem[155] = 144'h16891577e6a3e4d003beeb87fab8f1791185;
mem[156] = 144'h1449fbc8fe8d1f0118cffc65e80517e2eb9d;
mem[157] = 144'hfb601cce17f2fbf204c2e92ef660f15b10cd;
mem[158] = 144'hfe0b19dc1154e60101fff08611edfea9e130;
mem[159] = 144'h033c12cd10a61a1be0fff42c103be83dead4;
mem[160] = 144'h11f811a0e0bc05ff12b0e2911869e6221876;
mem[161] = 144'h046918eaf21311b9f6a81a78e58b0b37e92f;
mem[162] = 144'h05a11eafe71b0a34e4d00f48f83d0e1ff247;
mem[163] = 144'h1624fe58ef4dfe27010905b8f5a2eb2904f9;
mem[164] = 144'h18a6fbab1323e81cf2acf314ea16ef390bdc;
mem[165] = 144'h0ce70ca6f7e6e908faeef83c153414e5ed89;
mem[166] = 144'h1bf608d11405e5411a29fda706750670f828;
mem[167] = 144'heb8e0d36f9dbe922e36c13e6e2480cd219c7;
mem[168] = 144'hec7ff7381fc60b96f579fccf1bc609c0f326;
mem[169] = 144'hee6d16b8e08503cef6c30d48e93af482ed22;
mem[170] = 144'h13a3f085e91bf048e0a71d9dffd2fe74ff6a;
mem[171] = 144'h0b24198d1cb800ccfdfd113fea55108c1e83;
mem[172] = 144'hf0921805ecdf0e510e8af7310f5d0dc3059e;
mem[173] = 144'he66b15440433f5cf0b6e09041dee15d20c33;
mem[174] = 144'hf308e5eb1d3217eaf0d6002e0731ed7d1981;
mem[175] = 144'h1d37e786ee36186b1dec0c6c1ad7fef11eaf;
mem[176] = 144'he5df19e719c30908f65902381f02e4191c96;
mem[177] = 144'h1b1ae9641402ef5a1a5deb6bfe6fe1441b11;
mem[178] = 144'h07d8028406edfcf305b4e3951b3918cf05ff;
mem[179] = 144'h081de66a1213e33112fc02821f5b05531c00;
mem[180] = 144'h06180c25ed1f0529fe771fc8f28a04b1f9fd;
mem[181] = 144'he4b61930f4f202d5eda00ed0e3a4e9c603dd;
mem[182] = 144'hf7f904210452fc88e82114a2ed0800e805d2;
mem[183] = 144'hf7d7fa480c18e594fc64fd62fbea0c3be7c4;
mem[184] = 144'h1376eb94faa819b81a6af32709ba02570db3;
mem[185] = 144'h02670aa51611ed89f9eee5361c91e328f4b7;
mem[186] = 144'hfc4914fe0204f3a21a421f8ce73eeaa3f9c8;
mem[187] = 144'he4e20a59f2c3087cec85e619e1b20292e589;
mem[188] = 144'he01010320bce1f250e9808481e20f998e424;
mem[189] = 144'hf7b2fe0400e4e669ee4cebd51c3cee761b4d;
mem[190] = 144'hfa7b1a10fce60e6bfb62fdbceab30289ef60;
mem[191] = 144'hea5bf25bebff12e1fc88f0d508efebd81bf8;
mem[192] = 144'hf934e6b106f1fd5af940eed9198d0f171dce;
mem[193] = 144'h0f71e9ff1ff0f34f1439194303e7e67ae03a;
mem[194] = 144'h0fcf1a6418f202230b271075e3a6ea6cf7b7;
mem[195] = 144'h0664e3da179bffbd04e71bfce97fec3ae3f1;
mem[196] = 144'h0834006cff78ebcff90febc6ecb507a51fae;
mem[197] = 144'h1b8e0e7019d6179ff2071ae1038a066be6a2;
mem[198] = 144'hea56f6841bb7f39610a4fcc1f81515dcedd1;
mem[199] = 144'h005a1059fb371a0203f608061924179fe519;
mem[200] = 144'hf18b05ebe3741746e594029ceab218fcfa5d;
mem[201] = 144'h1816094814931d8afdf817b805a4ef5de183;
mem[202] = 144'hfb16f17a1aba145a0a38e47a0a7d03a3e026;
mem[203] = 144'h1f9511d6f3481ecc0f3ff8790dd4e7cf0624;
mem[204] = 144'h09e9f8a41d2c074a0801e486e3ede9040be9;
mem[205] = 144'he6290b3bf9a5e78af8cef7701832e27feea1;
mem[206] = 144'he0c205a708d4fd13051aea440e68e659ec00;
mem[207] = 144'hf10e033009b4ec2eeacbe595e97a0c18f3e8;
mem[208] = 144'h0888186803acfd37e53aeda2066af4f1f207;
mem[209] = 144'h0eb6fcb1ee3e1b9200bb017b020218741380;
mem[210] = 144'hf3cef4b3ff6201b5059ffda31f92ecd812eb;
mem[211] = 144'hed79172607eff141e443f056167af88d0a2d;
mem[212] = 144'h1d7b0de21667ffacf46903871ba3fd0a15a0;
mem[213] = 144'hf0150568fdd51c4e0bd5ffa5060715a6f2b5;
mem[214] = 144'he0eeedc1131bfcb7e5a81d4ae42ff2280b4b;
mem[215] = 144'h192d16e2ef4519d21dff1236f33ce1ff02a9;
mem[216] = 144'h08eaff351924098b034d07a5ef47e3791a6e;
mem[217] = 144'hf53805750d110427e8f1fa9809bfe4abeda2;
mem[218] = 144'h0f11111ce6f0e8c5f7d3eebd0486e339f4c8;
mem[219] = 144'h1187e01b001ae8bf0ad41cd60120e85c09e1;
mem[220] = 144'he6810e2a163deeade52c041607c8005811db;
mem[221] = 144'h1a43fba008fa045318d3f0caeb260f55fc67;
mem[222] = 144'h14d3f3c3167c04b41169194cec8cfcf0fb1b;
mem[223] = 144'heff3ee6d18c90bd5ea5bf9f211c10f68e1c0;
mem[224] = 144'h1dce0a7f1c081a611319188418ca0a62f1f1;
mem[225] = 144'he2daf68aff13fdcff7a8ed7af42306b90093;
mem[226] = 144'h1aa8f298f411084d0228e2e10aaf1872e4b5;
mem[227] = 144'hf040e489f5480bcaefe71a5d12611876e65d;
mem[228] = 144'hef58f347080bf578f99d05d8029b1048efbe;
mem[229] = 144'h0b0a1cf10086fd5410d1eb92f3a6f4a102d1;
mem[230] = 144'hf7721fc1f1b5f16e0bb2fcb31f3300100ab2;
mem[231] = 144'hf23715ab1190ef03e5c71b2ef59ae3df15fb;
mem[232] = 144'h0388efc219f8f9c116f9f2d5f8a9f2a008cc;
mem[233] = 144'hf7b8f4ef10f808eff718e222ea9e06921dcc;
mem[234] = 144'h1e2ae5ddee8e0ca5079cf1a4e9270b9bf71a;
mem[235] = 144'hf3f317ae177d034101b114edf112ffb80651;
mem[236] = 144'h0850f5d4e48deedefa80e0e40487f68a1f87;
mem[237] = 144'h1d1efe1e11cf001ee47def91f250ee200606;
mem[238] = 144'hf399005bec85e3def391ef5706ba1ddf1add;
mem[239] = 144'hf4ea0f610fe5ebe410efe54f17dc0bae10cf;
mem[240] = 144'h1bc5059700d90359fe991d2119f1eeb0e460;
mem[241] = 144'h135ceb3b15f9eed2fd6d1740f3bb0213e625;
mem[242] = 144'h1211184110c70961fe3f15e4077ffd911f89;
mem[243] = 144'h09ba1880f15c0fdf1a2803a8018ee01e06f4;
mem[244] = 144'hf45b0d2fedbfed3d182afff01cf70437faa8;
mem[245] = 144'hf020f70f12ddf0d6f6b8fe4cf76cf9fbeb93;
mem[246] = 144'hfb840d181fe6ef491a2fe46e010ce6d71050;
mem[247] = 144'h050b0b48eccc0080e11b1b61fff401a6e384;
mem[248] = 144'h043b1c56e7f8022bfa59f520f48604a3fc52;
mem[249] = 144'h1250eeef1115e075e7c0f8dd09a2ff49e74a;
mem[250] = 144'h0d920d211a5d1c27ea6c13d6e5101c4c0d53;
mem[251] = 144'hf073e4631e87ebae107e01c4fa7de190ede8;
mem[252] = 144'h145be79e04a2f70fe76cee84e33a04ccf57b;
mem[253] = 144'heaad19a3ea39f9ecf42d1fc7016017d90fc7;
mem[254] = 144'hf2141c430830e51ee8980bd317380e3f15ae;
mem[255] = 144'hf346e3bc1a7a19ae0811ecc1e926fc68e375;
mem[256] = 144'he17309a7143d0425e2c8f6d310d0f380e968;
mem[257] = 144'h0557f0c6e66fe53115b8f2b000790143097f;
mem[258] = 144'he67811dd1d15ec47f4b9ea8be977ebf411aa;
mem[259] = 144'hf50df935e20cf91118ee0f46e1350b88137b;
mem[260] = 144'hf2511a931e42e6bb1d01fd9bedeb11c9f7ae;
mem[261] = 144'h1c4de5b4e8a4ebca0641e4911f96fa87f1ab;
mem[262] = 144'hfb4c019e0e831d3ce9deec3c1c87f4fd1200;
mem[263] = 144'h1f7b0147f554033deec41f53f34ff749130d;
mem[264] = 144'h16d9ff15ed81e242fa3cdffb04f10015fd18;
mem[265] = 144'h0001051e1483ffcdfb4619ff1dea1890ef4f;
mem[266] = 144'hff1d16bae1b9f957e8fc1e6e003a0a621c41;
mem[267] = 144'h1bb004a6edece381efa008f6eab3ee41003d;
mem[268] = 144'h0b9cf27ef1d5e5a4e92dfb1c15c50ec7eeb0;
mem[269] = 144'hf7130bc10217e40ae53c1aab1d751fef0dfe;
mem[270] = 144'h03b21b411b87fab417a903dded20004c1015;
mem[271] = 144'h1d8906cee292e82ced21e1effc1efa441436;
mem[272] = 144'hf48f16c70952f2c90d00e5f30f00ea380e90;
mem[273] = 144'h0adfeac0fc99fcc3e67f1b831331109109a2;
mem[274] = 144'hf1f8f94d09001350fb95e759e1da0e56e076;
mem[275] = 144'h0179fc2917a303c31f530bc5f0dbf215e211;
mem[276] = 144'h1ac10d2c025ce9d5e048e9c709480efd12ad;
mem[277] = 144'hf405fe9ded2b0ca8eafc1a8b07a80506eee3;
mem[278] = 144'he108fa7ef25815c61c1803a8ede30a08076a;
mem[279] = 144'h1bcd1c13f61d08d9e3f51ab2ebd5020fe0c2;
mem[280] = 144'he67b1a310281e7c90a08e55b1f0a0e971811;
mem[281] = 144'he618107d0683f461ea3d007a1597ed1eee40;
mem[282] = 144'h16f9fa100cb0f814e839dfd201c7e75beffe;
mem[283] = 144'h04d505661fc211a31adbe692ef77f6b91f17;
mem[284] = 144'hf2d3f2afff78eabce7c612160edbfcdc1099;
mem[285] = 144'h054effc1f0f6e4de011a109410affaf709f9;
mem[286] = 144'h0fbb0955ec5c0c8c1923182dfe62e992f89b;
mem[287] = 144'hf813fb250b2f00f911d1eb8e04301934ebd0;
mem[288] = 144'hfc54e412ffebe9461b5c0f6d01adfc2e10e6;
mem[289] = 144'hf7b0ee67059efcfcecf01b381c000e51f63f;
mem[290] = 144'h1a151878ff0bec9510f4f16104a3188c18e4;
mem[291] = 144'he7fbf672efd90eddf4b6e8f11fe914920167;
mem[292] = 144'h13bfe885156b17e5067ef08c12521dc9e20e;
mem[293] = 144'h1bcfea7fec2ae7eeefe400c11445e83c0320;
mem[294] = 144'hf3afed6a05dc18751c411c9d0bf4181d13d6;
mem[295] = 144'h02ae0f92fc1904a80034fb8708d50cdef2e7;
mem[296] = 144'h180de8740082044cf4c01d1cf129fe34f83d;
mem[297] = 144'hf596ed47e5510af7f47f06c901f30b1809b8;
mem[298] = 144'hed841efbeaf2e3951d61fe341038e9e4054c;
mem[299] = 144'he56514760b4c0e87f2f60c7b107bea74e05c;
mem[300] = 144'h0d4514c2f8f2118a18b9f6d7137e1eb01774;
mem[301] = 144'heeaee22d1117e86cfa03095901b4efa1059e;
mem[302] = 144'h1cf7e58be963f7651ae0f5a11768f7edfc1f;
mem[303] = 144'h0eff0bbe1bb5093306761732f5f5035af837;
mem[304] = 144'h16a003451167f48cfdd9e2800d360b031de6;
mem[305] = 144'hf90c06dd19f11861f836f86beb5818040143;
mem[306] = 144'he722fb34fc2cfa531fc6f417e1e5131f1750;
mem[307] = 144'hfcfbe2121f1107251f351e540d7bf2d3f30d;
mem[308] = 144'h1e8f0a9714320e5c12470e3cf99e10d512f9;
mem[309] = 144'hf0eef08edfe2e9b0e35ef046064fe6ab03a7;
mem[310] = 144'hf175138a0ff11b4ffbee075dfddb10c6f291;
mem[311] = 144'h0eee0eb515ca0203eeb911a0097cf5b5ee11;
mem[312] = 144'h0eb9f3e5033d1f59e9a0ebed05131b730d3d;
mem[313] = 144'he3d0100f00d8e7ebf0430d8b02141d8a1c46;
mem[314] = 144'h0dbd0489055de8320710fe710f77f2ce10c2;
mem[315] = 144'h1ac80787f2680d24186ff28e15c3109dfea5;
mem[316] = 144'h0a8600291ac8fd15ebdbed77040711b10fcd;
mem[317] = 144'h1369f671180f14edf0601f560a13e48b1bd7;
mem[318] = 144'h12f71c50ea19fbaaf764e576ef05e3f20ead;
mem[319] = 144'he44e183d1c3811d4ec2815fe0ea805a5fcbe;
mem[320] = 144'h160c1c6e0a2707030a5ef73cf394e07b0b97;
mem[321] = 144'he98ee1890df31de4f0ede2681cb1f073f0ff;
mem[322] = 144'h1279fdc9ebe7ef16f0f406c80d8015ed0ca3;
mem[323] = 144'h1f840e6fe82a05330748fb27edf3f8f70a48;
mem[324] = 144'heb14f8090382e03b08dd1fc4158e0447e22e;
mem[325] = 144'h15d2e01516e50ceeeaa6f9e8e37ce92e07b6;
mem[326] = 144'h177df9d6fcd11d03efbc1413f05f13f5f0a7;
mem[327] = 144'h19a1e7dc13141ad21f0ffabfe1cc1e741eb9;
mem[328] = 144'hfc1bfa81e133f6f6fc5a0c8cf2a41d26e9fb;
mem[329] = 144'hf5f9fddd01f2e0dcf098f908fdef15ee1837;
mem[330] = 144'hf5d5f931174de687f47ce83aeb4d1b4b1dcc;
mem[331] = 144'h0a7d024c1b51f01e153ff98ffe851514064a;
mem[332] = 144'h1a5802400a80fbe6f286069019b7ed01002c;
mem[333] = 144'hf82cf7ee03cfe4a6e094e601f83dfb8708e1;
mem[334] = 144'he77bf39b035ef3ebf5ce0ee01c0609a1f0cb;
mem[335] = 144'h15f21f77e7721090033ce97c0f71ff7b01cc;
mem[336] = 144'h071d0c82facf0e0718aeeca5098f1833f829;
mem[337] = 144'h1e8e04da1dcef741e2940727ec3a1eb41df7;
mem[338] = 144'he68cfb32fc5cf16c12b10b5cedb3026f18a4;
mem[339] = 144'hf98df69f021ce48509bce4e009101cde0641;
mem[340] = 144'h13880028fb6d13dee77d038aea6f0661e12f;
mem[341] = 144'h099d10d7e0a4f9ac12d41d63e3cffc25e00b;
mem[342] = 144'h0df4e696e2a1e400e4930422158ffe9de3db;
mem[343] = 144'h1b9a05a20a9ce10506c30a7c05980993e5ee;
mem[344] = 144'hed3af9f110651aeb1e7e0b081ac50ae91ad0;
mem[345] = 144'h0d1b1f10029b020c01a2f2bc103005f6e80d;
mem[346] = 144'he9e10bc315431068f256f774f33913b70f71;
mem[347] = 144'hfdaa024ce1f0001a00abe2cdf26ce6c4ff10;
mem[348] = 144'h19910103faf1e115fdd3fbc10390f44704f0;
mem[349] = 144'h1988f217f25becb8fdb2ea890449f4b3ee51;
mem[350] = 144'h01aef5ff1b46e6c91af0e051f5e900140100;
mem[351] = 144'h12a7e7e8e575e1e8fddf0819fdb2f5f50f3d;
mem[352] = 144'he8d2e407f46a1937eb38e03ff68ae616fbdc;
mem[353] = 144'he514ef1411301ef3fc75062cffe10b27e673;
mem[354] = 144'h113bfd22ff3de08ee89d1f36f055ed6afdcd;
mem[355] = 144'he3f60907f83bf7f4067ce6e8e7c01575e3f0;
mem[356] = 144'hf752f989f2b5efb80d790932ed0305d8fca3;
mem[357] = 144'h08d210c8e086eff3e3ff0a0efbccfe33ec05;
mem[358] = 144'heeb717e41d2a1a1916a4026cf2a5f23b0e34;
mem[359] = 144'hf21bede8f037ed45fea0ec9f0a3d1c840e2f;
mem[360] = 144'hea021dd2fc35fde015b2f89ee75200d2e96c;
mem[361] = 144'h09c2f8b6f807fb8b0efc1f621b4d0658e471;
mem[362] = 144'h0cfbecbef814176de679ff03f28604d0e050;
mem[363] = 144'h00af1e50e600fa1ff4eceefc107ff6191a67;
mem[364] = 144'hf514eb901c90f9771419105808b5ed66f2b3;
mem[365] = 144'he99cfa3cf870fcd4e950120918a1f427ead6;
mem[366] = 144'h1c4cfa72e9f209611fd1f5bae51cea85e2c1;
mem[367] = 144'hf5d30883e431e98b1305fc31eca50f24fee2;
mem[368] = 144'hef47f4cc1966f3a413310b76099bf971f74a;
mem[369] = 144'hf180facfe4afe56009b9e7faff59e232e7d3;
mem[370] = 144'h0a5f0c82171d1b69e2461f921d5a01f3f7c8;
mem[371] = 144'hf2c011621229e226130f1e3903a118f91909;
mem[372] = 144'h03f61d78135f18b3e6420b92f6041d8c159a;
mem[373] = 144'hf361e10715c7f2d6e60a11400bff0bf3fe7b;
mem[374] = 144'hf415076bfeeb17970610e094e76efd05fc8c;
mem[375] = 144'h0f3ce23bf65b054c1325eb28e4a008ee1392;
mem[376] = 144'h0eb9ebe1f669fce7f13f1143fe5c134ff511;
mem[377] = 144'he93a1f1d12cb0ba5e693194119a2ff75e28e;
mem[378] = 144'h1b4cebae07c11fc80d171371123b0412f1ae;
mem[379] = 144'h1385e86cea9116c6fd1e0f080efbe08dee98;
mem[380] = 144'hf5850b2e13fe0c83f4bf006cfd58173500e1;
mem[381] = 144'h092bed75fd5e1f43ee4ff788003d0607f904;
mem[382] = 144'h0898f9abeb42130a1d64fc271697f9d8f5b5;
mem[383] = 144'h06891d68f6b1e2b5e8140b7906c8167ee65d;
mem[384] = 144'h15f2162ae9721a2e0382e510ece30bcbf67b;
mem[385] = 144'heb3f08db022ae55f1af61bbc19b1100c0c15;
mem[386] = 144'h1189e6450ddf014bfd10105febb11606e54f;
mem[387] = 144'h03590b561a81f9ff0716048a126f1bb01d03;
mem[388] = 144'hf275e7671f4815b7056d1cfbeff2fc4312f2;
mem[389] = 144'h0a11e7bd1125021bfbc8e7570b21f700e12a;
mem[390] = 144'h1eae07ebe553e0b504d7f28bf87df264e7ee;
mem[391] = 144'hf9882005fd200f72f7431d3718b2e3a8f60a;
mem[392] = 144'hf36e107418921d4ef13df0871337ee3ef5b0;
mem[393] = 144'he1f1016ff6321ec50f44e727f6760a74f66f;
mem[394] = 144'h123c1400f2ebe64e172d0ba5ef740364e793;
mem[395] = 144'h0e50049b01850e8b18360e24e43e07ddf4b2;
mem[396] = 144'h115b03011542122611941556ed911236e2cc;
mem[397] = 144'h032fe809ea420ab0e1d7e463fe260934fd56;
mem[398] = 144'h159e186c185a06afe678eb2512ad0f93ebae;
mem[399] = 144'h1e291454e6b01f8ae5770ed00484e627f13c;
mem[400] = 144'h0f81fcd004440357124ff59205c7e9d0eb9b;
mem[401] = 144'h000fe4d8168c1cb9f50ce3bc13f11445f634;
mem[402] = 144'h1b9d0ee007a6fdb40405f1961307edc81fd2;
mem[403] = 144'h0f5eff18f71d0a1af81ffef3fa86e847eb93;
mem[404] = 144'h0dff03eb0089f6c2163ef773f6200c521bf6;
mem[405] = 144'h1e61e55716dbea77e0bdf0d9f6f8f3cffe65;
mem[406] = 144'h1c55f302e368ef6bf68009e8ed9ef6df0d58;
mem[407] = 144'h1208f8160d2d01ac09971ec80d46fb3d1d81;
mem[408] = 144'h041e1c981d6e082701e8ed5e14ce189d1ab6;
mem[409] = 144'hebee0e0a00f9f5930603192116a6f8ca0ff2;
mem[410] = 144'h195f0c67fec8eb0ae0a9e156031b1c27e87c;
mem[411] = 144'h0830fb6b03a0f64af4810bf31f5eedc4e354;
mem[412] = 144'h1972ea90e0f30bf902b8e1bb200dee0ef92a;
mem[413] = 144'h0fa7f7e5076cfce21c53f924fdace242161b;
mem[414] = 144'hf973f523e71de0e5f7e1fcbe04f8fa0c12f2;
mem[415] = 144'h19b818daf040ea8aeb1f1602056307dc1735;
mem[416] = 144'h1f1fe5aefc81e7ad1e2df0fffcbb11d61513;
mem[417] = 144'he8c4e06402d30d350903067a0e20184ee0fa;
mem[418] = 144'heb52e852e5bf0182eec71d0fe2900ddf17ab;
mem[419] = 144'hf46113fa1a4f04d1eb2d0948e55bf64ae4b5;
mem[420] = 144'hf506fde7ec36f42deec4fe081f21ef18ece2;
mem[421] = 144'h0ce2e4ff1bbee13aeb0113ecff72e2a2e4e7;
mem[422] = 144'h11790bc608601b85175617cc008c073d1ed8;
mem[423] = 144'he15e1d6dfff11d4ce4a51c40009ffe421267;
mem[424] = 144'h038c0466052016b50c5e126ff7ee0df7ef82;
mem[425] = 144'h0021f090f3aef885f06408940fd4f0731d20;
mem[426] = 144'hf6c2e53c011dff020b42e888edf40a25f865;
mem[427] = 144'h1800e4931f7507a2ebc1f5b6e28ae857042d;
mem[428] = 144'h0b47e3e100c9195216c811e4f08af2aa174c;
mem[429] = 144'h15a41a25faa5e40df55fe2ae12720c040221;
mem[430] = 144'hf67f01c901befab6074012f1ea2f14f217bd;
mem[431] = 144'heff4f9fd1a2be20bf32413cce213111bffa2;
mem[432] = 144'h096605c30d10e2eee7e312bef43ae7e01511;
mem[433] = 144'h0f16ec58e4550af30d21fb7f04ebe488eef5;
mem[434] = 144'he14effbee727f58ee944fa4ff3c81731e001;
mem[435] = 144'hff9be4dde7a01e76e3d5edf605930dac1f3c;
mem[436] = 144'h0b54ea2c02a2e9deec8be83a07ef11521736;
mem[437] = 144'hf66805c2e0f7e0141ecf1089eb0f1ca4f00b;
mem[438] = 144'h1531fb30f383fd73e4560da00148fa88fc1b;
mem[439] = 144'he546fb16f64c1f19e7fbf333143a1d2bfda6;
mem[440] = 144'h0d7ee51000c4f566fade16e9f29b14d81136;
mem[441] = 144'hed2c1db21ff10fc9e48c1c94ee5c010ef9b7;
mem[442] = 144'he23a0a64ea341bfceaf008b90a7af4ae0e25;
mem[443] = 144'h08a5f29af8e9f35c0bb3ffcb11ae17581666;
mem[444] = 144'hf33de8f4e24bf9fc1ba8f4f9ee3b1823143a;
mem[445] = 144'h1cad122c13a70859170e1671fd87fa1be490;
mem[446] = 144'hed1de913fb2a1deb109ce5a00ed31b8a1abb;
mem[447] = 144'hee41f7c9e8fb03170dbffa85eba0ff3f1272;
mem[448] = 144'he984fdba1bece2b8e5b0ee500b86f28df66d;
mem[449] = 144'hf180f63ee0b8fea71f141368fa0f0bef091f;
mem[450] = 144'h155af09e04d6f5460b55eddd1de4fe290b85;
mem[451] = 144'h083ce1d0e23bfc44e9c00c7908ea0802fb63;
mem[452] = 144'h1559019defebf8dce26ce51c0629ea3df05f;
mem[453] = 144'h0f1bffbeec26000902c9fb15e72ae4c60532;
mem[454] = 144'he3910ec70f60fca8ecde0efa1ad11af8eafd;
mem[455] = 144'hef65ea87139d1319eb5c1b48e39e0492fa65;
mem[456] = 144'h1f1fe3f0f42702f106b3f330f7f8e71ce7e3;
mem[457] = 144'h15541b4b02dd0e010786fb9115e6feb60cd3;
mem[458] = 144'h16c100b0ff2c009d0471fa90117be25104c5;
mem[459] = 144'hf2ef1ac8f4bc0916173fefda1e49ec170fdc;
mem[460] = 144'he1d31dd7fd7fff28f628feb21bb4f6a009be;
mem[461] = 144'hef53f9b3067febdddffff34dfa3907d4f6a2;
mem[462] = 144'h1caa1b55ea01f58b0841fa82089a0233f0a8;
mem[463] = 144'h10f702881451f4770431e89f0434fcccf249;
mem[464] = 144'h1281feb41cc4e26f05110ec0ea8e09b9e2d4;
mem[465] = 144'heded156604e9e8f9008410d6fd0bfc7b0f45;
mem[466] = 144'hfe4c05e4fd8a1f40f6ab0840f11afd7c09e7;
mem[467] = 144'h1034fbbf19e411c8f88befbbe803155a1093;
mem[468] = 144'he2b8f477f90ff38c14f702d104f2e509e3d2;
mem[469] = 144'hf2b5ff3c0c2d1ab91a990c2304b91cc6e9aa;
mem[470] = 144'he91c087f0407e4941a2010401c7ef48de082;
mem[471] = 144'hf1e2f0b7eb0e0e8cf30601c9f0f0e246e0b3;
mem[472] = 144'hff040844f4c107ef067314b11f2103fd099f;
mem[473] = 144'h0b11ea50002e1efde483fb61ee5e1d7000df;
mem[474] = 144'hf5c9eab615d4edd81069e4b21d0f1e311a85;
mem[475] = 144'heb10e685e9c5f650023a050ffa8ae6bdfee0;
mem[476] = 144'heaac0322f85c1a7802940d5bf4c51bafef9d;
mem[477] = 144'h0f16f02f0973e3e9f0aa05af15cbf2321b50;
mem[478] = 144'h17020ee9f900fcf81a65051f127ffb6a1e72;
mem[479] = 144'h1f1905960931181def9fe885e993efc01b1c;
mem[480] = 144'hfa2c0060f0adf1bc185d05960d0f1c3e01db;
mem[481] = 144'hfb5df92703b60eadf28f17e5fcaeebcde43d;
mem[482] = 144'he6b5ee8e02e3fe5100aae0f1e7cd1c4dfa5a;
mem[483] = 144'h0c66e92e1b910470e0d0088a175fee1c1b15;
mem[484] = 144'h1db51202ed39148ee1cf0b07f9cbf3e21dff;
mem[485] = 144'hfe2209441e6e1c891e4d0c36f819eee0fa41;
mem[486] = 144'h00481a8c0d99002eec53e4011cd11010f1be;
mem[487] = 144'hf1c3f3ddedc4e9fa147b16e8ef4f135bf871;
mem[488] = 144'h0f9eeca8e49d143516260005fbb217eaf794;
mem[489] = 144'he0f5e490e458fbe5e7fe18a3103ee56b00a7;
mem[490] = 144'h0f33e32f0a74e349ea29178112b9fdae0ac4;
mem[491] = 144'hf7a60792e9e3e53fe363ee11f3f2ff84fe3c;
mem[492] = 144'h1d9a05fe08210481172a13f41857137f1fb4;
mem[493] = 144'hf0cce1dd1ace1139e204f256f898f69efa7e;
mem[494] = 144'hfc541742f10be775e2271a120918ecc2e8f8;
mem[495] = 144'h00781a6cf3a4ec7bfaea03d80f75170510df;
mem[496] = 144'hfa7eecaef08a1cdcfbdd13f119e40a4e1f61;
mem[497] = 144'hf00903a200f3e0b6ebf21ccd0e5c09a5f603;
mem[498] = 144'he5b21d20e26f0fcc0c76e2c506df0836fe7d;
mem[499] = 144'he8c313b705c2e1591dc91d73ff38f47017d1;
mem[500] = 144'he876e407124af1eaf78115fc02e9f4c0e431;
mem[501] = 144'h108415ce04d1f5f9e7d6ebb3f6e0e5781927;
mem[502] = 144'h0b27f1030953f85fe86411d2ffc6ed25fc9f;
mem[503] = 144'hf4e9ec74161b16550bfff179129df591e2df;
mem[504] = 144'h021d1021fbcffb52f15ff566142f144d1d96;
mem[505] = 144'hfedced0ffbf8037c133f1894f9c5ed21e5f3;
mem[506] = 144'hfd44f974f94e0999fff2f69af68b05d3fbe6;
mem[507] = 144'hf8c6fd98f6eb0203e07a03ab06a60ebff1b4;
mem[508] = 144'hfb8d0003fd7c0dfde5cf1ab7f4e416eaffa9;
mem[509] = 144'heb4117ef0dc5ed8c1267f3c5184b08bef79d;
mem[510] = 144'hebc41ed6f0aae2b6168ce0a814e805cde8e0;
mem[511] = 144'h0549f42b17c9f2ac1138e31d0037e83401f7;
mem[512] = 144'hef19fda5f4e8009905c2f719fe9b0a70e697;
mem[513] = 144'hf8e8e648f7d4154b126fe9cbea96f41618b2;
mem[514] = 144'he756e3e505150ae00617eb860943138bf8d9;
mem[515] = 144'h1a0be01be39d00c7f45a0e76f1a9ee0a1da8;
mem[516] = 144'he8c207d4fe48167eeb30064b11c1eb52eeb1;
mem[517] = 144'h0263e10303fd02b5e056e0c0e6090e9f16af;
mem[518] = 144'heb3ae086f3a3f6581199e10e04e4f36fe295;
mem[519] = 144'h0c08e787fbb8e3401c811c24ec2df3d915ec;
mem[520] = 144'h1ef3f4f805fee2e4f86fe94be3fee46af841;
mem[521] = 144'he6fc02b9eb0b19b6fee4ffc3f5baebdf0683;
mem[522] = 144'he945e497e8a5f9c4e469175409430e1a1f3f;
mem[523] = 144'h03fb1dc20d7e095deedef0a7e87b17aa0455;
mem[524] = 144'h1207f51ceeb4090fe45de046fc8601ca08e1;
mem[525] = 144'hfc4408dd0e8a0b4e027e04060f41ffd51673;
mem[526] = 144'h054fe8e9ebed1fd8e0871135e282fcbdfddb;
mem[527] = 144'h1672f39bf2c0071712d20f20e8b11ff00ba0;
mem[528] = 144'hfc30092402b414931a9ee8f0e05b0d051530;
mem[529] = 144'h0943e8d106dc1914fbf0f84e1342ed950134;
mem[530] = 144'heabfebb7083e12eb0064ecd417f6f9b1fcee;
mem[531] = 144'hf83fe6281875fa151d271e0ef3eee1cbf2fe;
mem[532] = 144'h09c108c5fe45ec7f0043e3fefe1befbfe21e;
mem[533] = 144'h13f816061c45f65fe0e8e1d91f1a104102bc;
mem[534] = 144'hf8f90e9502cae06b0dacf65e1f5ef132e3a7;
mem[535] = 144'hf4311c7e1c2909390ecd0151168b0154e3e0;
mem[536] = 144'he7cffd63f61c12be16e3f0d0fb5a02fa059f;
mem[537] = 144'head2fdfae2dae772e388f43be9a014d7e0ae;
mem[538] = 144'h11b70561f992ee21e7e9f545e3f2e0bfeeee;
mem[539] = 144'h07b51f56ee57f7beed70e296ebadf7691321;
mem[540] = 144'hfc7b1e2cf2ce05ce1fe011470065f45e1593;
mem[541] = 144'h0f481c26f06d117ff79aee49102d0408130b;
mem[542] = 144'hfe9e1847fa3b04e0e2cd088011a6e52f0839;
mem[543] = 144'h013b06e5f052ea260128ffc1ed27013ce8b6;
mem[544] = 144'hf6491564f5451293eaa10bfff57607df1833;
mem[545] = 144'h01911bb7e335e93fe39c1f4611cd0888f4b4;
mem[546] = 144'h1e3e07f4fed8f17111b10e0a196ef492e1b6;
mem[547] = 144'h01e5fafd165eee12e1da10c70aa90b890d71;
mem[548] = 144'hf521e5310df7f6b8ffbe0f36e5a81f7ae82e;
mem[549] = 144'he99e11460bed00331e48e67ffb101947fd78;
mem[550] = 144'h1ac013d3130a1143fe050abf046a0c5ce2cf;
mem[551] = 144'h195dfc261213fc48e298fed01fe80538eb13;
mem[552] = 144'h1cdcfd69ffcf122aed450996e1431f2dfb35;
mem[553] = 144'hea57f22febeee4ef0aadf5c3f02df37e193e;
mem[554] = 144'hf432e54ced83e3130a320c82e63b1522ee82;
mem[555] = 144'h0b69152de8c8062ef0d2e523fd1704cd00d3;
mem[556] = 144'h0dc30b1418710f8308d6053a025c1587eedc;
mem[557] = 144'h1836113be9a41090e2f90ac201ac0ed3f66a;
mem[558] = 144'hf8f41a3210d4fab8eccd1070152af717f704;
mem[559] = 144'he27210ed066103c801cef57c1b490bd6163e;
mem[560] = 144'h0be100f0180e09611b35fdcef678e9df12b8;
mem[561] = 144'h13800a570087e6f81ac1f52b0b73e2b0012a;
mem[562] = 144'hf24ef2a6ea47f22c0bdafc58e367f83ffb38;
mem[563] = 144'h1f46ef0c0466eec0f96c019b0002f25019ac;
mem[564] = 144'h1e92162ae831f624175ae9d41bc507200b86;
mem[565] = 144'hecdef283f532e5bcf70e15f510ff0697e990;
mem[566] = 144'h1d97f81a0b661e21f6dd0549074ceaae09f2;
mem[567] = 144'h07141fd11500e0db1c7ef13f03eb09071f48;
mem[568] = 144'he879f567fa450b77e8cee50cf86c1280e1e3;
mem[569] = 144'hf6991a0ef95a15eee375ffa713e503a4e39b;
mem[570] = 144'he6fe0c48f44efddbff0b094d0bf50828facd;
mem[571] = 144'hf92cffe50fc2fbfce715157ef4cef0031fb6;
mem[572] = 144'hea48e713eddb120011f3f4ef00b7e08315b2;
mem[573] = 144'he4f80c7de0331a5300a306beff4ef66d11b1;
mem[574] = 144'h00d3f2860c6c132e14fd0e03f6e8f0ab1bd0;
mem[575] = 144'h1995ede707d0f55bf391eb78e30404cff6ae;
mem[576] = 144'he99b05d80575ea0d043a01fe094f0f2a12e4;
mem[577] = 144'h1243e497f66ae1d0e69c0141fb84162aeba7;
mem[578] = 144'h0655e8c810480de8f473161d109c0e04e6c6;
mem[579] = 144'h1d531d34fd7afc11f1c8fc98fc6de1f917f3;
mem[580] = 144'h0a74172a1cda057b048ee572e2cafeeae1d0;
mem[581] = 144'h10eb0cdcf5c4f1bdfc71e6a00fb3fed4ff4a;
mem[582] = 144'h10a5f4751e54f765e8a512cbe99a0205e203;
mem[583] = 144'hed26fa8ef19fe97a1c6e07def7d60360f5e4;
mem[584] = 144'he7c00c5ff1cd1cd8177913e9fa81ef21f11c;
mem[585] = 144'hfcbef61de9f2f4ac1316e981f1761900ec08;
mem[586] = 144'h1f05e6fa15520482ffd103f51ab61fcdec8d;
mem[587] = 144'h1a3a16551b3debbcef52f83ffe86184f0b6c;
mem[588] = 144'h08880dcf018aedddf5d8f41ae43c1093e84c;
mem[589] = 144'h04b1e633056a19b619ab12b2e9210ba9e31a;
mem[590] = 144'h06fe0404ed9ef703f7950b78e9c6f8d50c98;
mem[591] = 144'h037bfce513e0e9510f51092cf7b4f3f20f5d;
mem[592] = 144'hf9b60610f3a8fa2405f503b9189a0d72faf4;
mem[593] = 144'h1ade1915e99ceed80a72e7b3f7a807200af7;
mem[594] = 144'h1693ec0f12e4ebd11546f9031703ec77e2c4;
mem[595] = 144'h1459f7c8e4541ae3f72f08e4f4d9f2351508;
mem[596] = 144'h1a9a108f0f08fd33eaf2e3230984efa21686;
mem[597] = 144'hf39e1aaf1ba7f83afba1f48a176cf48b046d;
mem[598] = 144'he4ed192d0a41fbd6e72fe523f3a8ece2171e;
mem[599] = 144'h1c9e0149f8d9079ae6001d331ff9e1a6022c;
mem[600] = 144'h1a88084615fdf94011b2059403fff903f665;
mem[601] = 144'h158e02ed0b0dfdeb0843e2e6eb2a1839ef06;
mem[602] = 144'hf4c7e54202b20eb5f72c1b8ef9e1e397e8d8;
mem[603] = 144'h050b187c1fa9f6e8f96eff4fe33fe2e1fb7a;
mem[604] = 144'he4b7197919d91db3005c0c2a06dcf6ee0b89;
mem[605] = 144'hf4700fe2031e05a20521e34b1e1c1e8405c1;
mem[606] = 144'h0a2ffdaee5d2048efda6ffb2e1df003e0cca;
mem[607] = 144'he158167de4e80bbcf065057ae1ccfbc2eedb;
mem[608] = 144'he097109ef6330d250e130831f1be10ca088f;
mem[609] = 144'hf25f14890762174bee6f128c1a840064e347;
mem[610] = 144'hefb81d34f29a155b0a4b1596fedfff480397;
mem[611] = 144'hfb21ff71f886f46911f1f3a60437e73ee241;
mem[612] = 144'he93a1c040798e2761a22e5250eea1e55f210;
mem[613] = 144'hff351bc7f3ab1236ed210eb113c5fda5f5da;
mem[614] = 144'hfad2fdeeefc817bcfee3e4db0e79ea0fec8d;
mem[615] = 144'h04dde9521bbf1bafe85dfc0208a1fbc91c35;
mem[616] = 144'h1c9ce758e340e82510ba0fe3185ae8231526;
mem[617] = 144'h1acae472eb8a0d8bfa5318731e44f9dfe422;
mem[618] = 144'h1ef01c37ea361e18e95b0594eb59f498f078;
mem[619] = 144'h0547001304bc1b4111ba184de1570631039c;
mem[620] = 144'hfffa1ea516c9ee35f8cce8f206d905b61e3d;
mem[621] = 144'h12f9e601f7cefc8cdf9fe7781862f37eea1f;
mem[622] = 144'hf4731c08fab31c97e33a0fd1e63f12981657;
mem[623] = 144'h1bb10727e691ee7617461f7b0313e1c7e9a1;
mem[624] = 144'h0fee0ef2f869fc951a0119320bb20c0e1d6e;
mem[625] = 144'h03c10ed71f0ef32e00bf157a079a154ef250;
mem[626] = 144'h0ecaf3190080eadc05940fd0e4d9e7bc0720;
mem[627] = 144'h145bf11f0f63f235fc8cfc65e0fae49619fe;
mem[628] = 144'he6a9097303f2f8520a79eda7e5f70dc9fb02;
mem[629] = 144'h0863f102e28de957fe1df743013cfd47fabf;
mem[630] = 144'heb221b01fcdae5cd1b45fff9041b1072eec9;
mem[631] = 144'he984fd1afc8908e9f7821825fce7ee22e275;
mem[632] = 144'h0ae8e3bd0ee709ce061b09baff24e6b7f81f;
mem[633] = 144'h117efc9417c3fd00e91ae57f0b4ee414e9cd;
mem[634] = 144'hec49ff22e88e002f0caefa13e4231f0df25a;
mem[635] = 144'h1fd902080911e91503521e53e563ef8def87;
mem[636] = 144'h166915871c5f04e314e0f548f83bff4cf8a1;
mem[637] = 144'hf800f3431d3815d7e27f0684028be2b91c08;
mem[638] = 144'hfffce19f177904b6f4f611adf38ff95cf0fb;
mem[639] = 144'h0c05fe7f1be50d87146a0c3819111260e3f7;
mem[640] = 144'hfd3806f21ed6f01c18e9e5a5023cff0a0105;
mem[641] = 144'hf4aced01edf717f4e9b9ed63f6a50fd91444;
mem[642] = 144'hf99eef39ef1d1d02e138055be5cae8e60f47;
mem[643] = 144'hfc7104e1016ef748e3a70a8c0360052f0830;
mem[644] = 144'h1c241fbfee9402fa002cf8de12460cb209d0;
mem[645] = 144'hfaa1e9b40495f9230c390093f06805bceb50;
mem[646] = 144'hf0990b07f0201d5cee77eb31e9531a8be5ff;
mem[647] = 144'hf4f41d36f0d71adee88f0cc60f6d0c4eeb24;
mem[648] = 144'h03e6fb8a1cd41909f4371e1210c7f5321b93;
mem[649] = 144'he1bb0bde1123f4050793eb9ae392162af898;
mem[650] = 144'hf30ee19b1057f7eae0c5012fe46211d9fa5e;
mem[651] = 144'h1ed0ea4c03be1f60fe1f13900ee216dbf4fd;
mem[652] = 144'hdfde10dde9f80346f8681dc30293e62be0b4;
mem[653] = 144'he1f1e41207c71b8bf2db03ff1af1fb1aed5f;
mem[654] = 144'h1b6a1604e468e475e602edeb1e1e1e5aec9b;
mem[655] = 144'h06faf2860920f8c4041e0f5e1a9af1c50f84;
mem[656] = 144'hfa06034df5cae2dbe8ad0f35e2b4fc76e90d;
mem[657] = 144'h041a03c2014b0a16efb20d0cf9461f6b037b;
mem[658] = 144'hf3e10a37ec530e3e1591ea44eccf1c9bf071;
mem[659] = 144'hf8560149ffcbfff5e31314a11be5e0b404a5;
mem[660] = 144'h0f020f1e18a5e45e149df26e1b30eb311afb;
mem[661] = 144'hec40f77c09991b68fc91f092187e0f02156d;
mem[662] = 144'hfa9be7fb10ac0187e5bae5a8034dee101a98;
mem[663] = 144'hf66ce1770f2c0f69000afe82efc00958eadf;
mem[664] = 144'he9fe1ba0f4bfea5008981e8a0ae10fb00236;
mem[665] = 144'h1b2ae403fde5e16415060aabfe53eefbeb8a;
mem[666] = 144'h1e1007ef08a91053eacf183119d00e21ed1f;
mem[667] = 144'h03e0099c198dec73e92e018b135511b21596;
mem[668] = 144'h07d6e961f8f409ac1b18f6e8fa46e2f5069e;
mem[669] = 144'h1d99f4540c9f1a6319e6f6e80ed6f54ffa1b;
mem[670] = 144'he956e15ae618e9effbd906e11723f65ae7cb;
mem[671] = 144'hedb4ebcb0126f3610caf19bde953f7ff1beb;
mem[672] = 144'hf550f1490c821d5aefbc18cef37e0fe3f0f1;
mem[673] = 144'h1496ed5d11f8036feb55fc34114fe453f773;
mem[674] = 144'h09d8e04613c2e898e74c01d911d008610e7b;
mem[675] = 144'h0d431ea61522141101f9f46bfed515fc0f3e;
mem[676] = 144'he17de3ae00e6eda6f26ae995041dfe1bf2b6;
mem[677] = 144'he462ee430f47efeefab804ef16441ff50b40;
mem[678] = 144'heee3fd29016cf4f90074ed960804eaccea6c;
mem[679] = 144'h0497e013038ef83c0dd5f8ec1400fad611bd;
mem[680] = 144'h0c96e6d51767020a0fe90ce013c2fa620ded;
mem[681] = 144'h04a20472fae8e05be706f3dde47be39fe257;
mem[682] = 144'h1926efc30cbffb59eaa2fd84fb490f1bf5bb;
mem[683] = 144'h10ddece2e150f930f31a15f0ecbef8851155;
mem[684] = 144'he41ee36e1fe90f14f91117c8e088feca0a0c;
mem[685] = 144'h1a2c1401fde2f908ebf810fcfb16feb503e2;
mem[686] = 144'h11890045fb4110e71b5a11c6e347f65f006d;
mem[687] = 144'he4b2e9f30efbee6c1ddef28d0850f191fa67;
mem[688] = 144'hf987f59d1d8f0e9cf769e0b9f4ea130ee4f8;
mem[689] = 144'h1b2ce359e8b41a2ce4bef26e0b2ae356ecc2;
mem[690] = 144'hf8fbe4f5e441169915c7fd97fa0afc0c0da4;
mem[691] = 144'hef480a49e112ef0511100a0af505e43a0087;
mem[692] = 144'he6ebe099facb116718620890fd1213871de0;
mem[693] = 144'he6d6e1581d2a0ed7eebafdffe16114faebde;
mem[694] = 144'heae2f594e6f4ff6cf342035a0bbe1326f69f;
mem[695] = 144'h0c0b01c5007ef71c07d5f906fd4718bde22d;
mem[696] = 144'hfa25e135f459fdb91848e7bb1f6f16d2fa74;
mem[697] = 144'h191cfc921a70e4450fa316bcf89015a2ea94;
mem[698] = 144'h0a48f86e1e43079a1b33fbcdfa85e6d40038;
mem[699] = 144'hf03c1c3bf6e9f938e40c087d1aa903d91bfe;
mem[700] = 144'h1aef01f6eb9ff6c9062c05d9085c1c8ae023;
mem[701] = 144'h1bd6116a1fc215a4f86c052fe0d81611fa65;
mem[702] = 144'h063dea33eb20e2dd0fbeff20f80412c8e07f;
mem[703] = 144'h1be9060310c5f7afea430c3418eb15be1e7d;
mem[704] = 144'hf91913aaf23d1361f5fa12521d431f0eecce;
mem[705] = 144'hea0df3a31d9a001b1323040d013313e60c64;
mem[706] = 144'he79cf3c4ec7d1ba1f599f84a14ed0d42003d;
mem[707] = 144'heb3f1629f0e6e16d075400531365fefb1759;
mem[708] = 144'he6df152e119f08580203e74712c9e70511e2;
mem[709] = 144'hfba5eb6bf396f3a1170f0ec6e3d7f1e4071d;
mem[710] = 144'hfbd113860bec0d631198e5ad0b1c0721e536;
mem[711] = 144'hfd161234f6301b4de6dfea7b0f1a04bfff62;
mem[712] = 144'h05370b8eef84f1c2f884140e14fe05caff55;
mem[713] = 144'h1880e0f1f373e2eeedb00e4307b8e61fe50f;
mem[714] = 144'h09a5f2f0fa7615680d4e05e9029618051aee;
mem[715] = 144'hff531f5de94de3d6127503271953e5991957;
mem[716] = 144'h14e11049fb52fdedf3cd087c0ed112a305a0;
mem[717] = 144'h121e0e86fe28f9cafdabed85f5dfeb75f137;
mem[718] = 144'hf6fbf4ad078c0fd1fe2b1c68ebc0e4edeeba;
mem[719] = 144'h110ce1e9ff63fd1d0ae811ccf3f9e354f5a5;
mem[720] = 144'h1e44f2100198fe2e16b9f12e02cdfa9600f2;
mem[721] = 144'he8f7fab714c91ddef93c058d07131266f347;
mem[722] = 144'h1eaaee621e8a041cfb7fe5fbe98001f21924;
mem[723] = 144'hef42e594e915f3481bb3ea1be932ea65e8fa;
mem[724] = 144'hf209f5710c9f13c2e5ed0f02f22912e1e586;
mem[725] = 144'hf965efdf108ffe441c2ae6b30c03153e0d21;
mem[726] = 144'hee7501ad0a67ec39e07ce4e1f2d01181062e;
mem[727] = 144'hf318f01be04efa21f782f8be0366f0130fcf;
mem[728] = 144'h1f6f0f33ef23137fe6720f00ed640b7603d5;
mem[729] = 144'h112611abfe2100180c6ee3da19dfebd3145b;
mem[730] = 144'hf714e97aef0de67aea4ae4d9141b178d1b2e;
mem[731] = 144'he4581a5afbb5f005f4afffe8057905d11aa1;
mem[732] = 144'h1528e7e8f0b61f4bf0fdf40612bd06a6ea65;
mem[733] = 144'h12b409df1f6be1340c971fe6eb99f0a31100;
mem[734] = 144'hfd6dfab2eb18e30aeef704be1111ef56e1c6;
mem[735] = 144'heaa8ff91e0dd11fd0a3dfbb8f9fc04bcf716;
mem[736] = 144'hfdcc0986efc812bd0d131ef2e96900f70d3b;
mem[737] = 144'h04e4f8c11b83fba1e96c00bcf4351135fa37;
mem[738] = 144'h012b0c7f04cef98612cdf0960ee809c111e1;
mem[739] = 144'hf226fb10e21cf3131205f386e508fb010a0e;
mem[740] = 144'h1738f1371f61e160fef218f61f7f178eeb73;
mem[741] = 144'hf0191fb2f1ff0a24f43f1eb4f0af01cee1d0;
mem[742] = 144'h1c99e63f19f80400f0131c27e9190373f8b9;
mem[743] = 144'h10571aa0f218e108e64eefac044cfc0f1112;
mem[744] = 144'he114ef84f6c3fb230f941ba41803023e020d;
mem[745] = 144'heb5d03721603ef9e09480f2e11f1e412eba7;
mem[746] = 144'h0c8be85fea4a0051f48ee24aff80e3ebfb77;
mem[747] = 144'he8fb00a308f50060fe35fac90b94f85416c3;
mem[748] = 144'h10c3f640f4d9fb431898e8cffd721731e742;
mem[749] = 144'hf954198d1c3dfaa2efbcf4c7f613e0b8ed36;
mem[750] = 144'h070415260f16ec22fb91e20fe0cef2f2efa7;
mem[751] = 144'heaf2e3681434e1ebf0810635e7a3fc3be40e;
mem[752] = 144'heec3ffe8f1b8e6250a9b1243f6520a7f0fdd;
mem[753] = 144'h0ede1833032bf442179e0ba8f273f20ded7f;
mem[754] = 144'h007f0cd10553fc43e90ff57ee99811ceffac;
mem[755] = 144'he29ae2a6f28414dc1050e6bafc82173c05f4;
mem[756] = 144'he706e6ee05f2e0c1f498fc591f1ae63bec2e;
mem[757] = 144'h091709ea19b90bc21e1efa96e157e07a0156;
mem[758] = 144'hf829fd17ff5907880a9300851da7f2cbfe27;
mem[759] = 144'h1f0005071619e5a2141813e018d7f9a6f39d;
mem[760] = 144'h07cc186debcce476eaefe63ee87ce5e80007;
mem[761] = 144'hfd68e137ebaaf733eccd0c70052104041642;
mem[762] = 144'h015be44ee8c2142c0c35f2d2f979119efa38;
mem[763] = 144'h15edf5e4e01de57f0c691fce156de3901ea2;
mem[764] = 144'h0ca30f6fe6af0d370149086df1611f7ce792;
mem[765] = 144'hee6fe859e8c204ae157a07af0bfa097d0756;
mem[766] = 144'hfc1215031edc1ab906ce0dc5135c1f4f07e0;
mem[767] = 144'hfc97ec741dc8153d020b0b4de426fe1917d6;
mem[768] = 144'hf514e41a076cfab0018c0b61f65816df1896;
mem[769] = 144'h02d21cc2fdfde62be7c4fe7913960626f207;
mem[770] = 144'hf4cd16841ccd0ce806ebf80215a9078e10bd;
mem[771] = 144'h034a06891935e8bbf4e117b8fdcb0a0300db;
mem[772] = 144'h04beeba0ea01f98602c2fa1e0251e437e659;
mem[773] = 144'h096ee78b0aebfbfd18d812df05df1073f095;
mem[774] = 144'hf6ff1d8ffda7e9bcec8c1eef048405cc1f26;
mem[775] = 144'hfce315cdf4260d2d1ff1f44deddeffa1ec9c;
mem[776] = 144'he90005ff041ee952110c10dcf8c6f908e2eb;
mem[777] = 144'h07d9f5d3f8461711029219e10be91825ef10;
mem[778] = 144'hf022135ce82bf854fced1071f608e6751fbd;
mem[779] = 144'h16fc157d0081148eeb8d1203104ffa47fe3c;
mem[780] = 144'h132c0442e59deeb2068e132deea8e8011218;
mem[781] = 144'he8ccf8b5f49eec25f9a60f02f5b60b681c38;
mem[782] = 144'he179ec50e0d3e12ffb420c3c1b6bfd2916bc;
mem[783] = 144'hf7970549eca0108a0fc318b30e8fe8850697;
mem[784] = 144'h085a0312066de562162c1a360a79e26a003c;
mem[785] = 144'h0bbdfecde608130e1b0016e9fa99e71e1578;
mem[786] = 144'heca003c8e667f0a51b8fe95c02e700220ab1;
mem[787] = 144'h1c520ed0ea70142201680b740f261d99efa8;
mem[788] = 144'h1b01f890e85fed6c1d3bfa7d193ee3dc1a3c;
mem[789] = 144'h07d414c9f2a9e181149dfb93e28916700087;
mem[790] = 144'h1f6ffca00a751cf71f970e06ed1dea7aea7b;
mem[791] = 144'hed97e0481c3f199008e003ed0733fa1e0016;
mem[792] = 144'h136f05a915f9018b0b88f877e8adfc9f15e4;
mem[793] = 144'hfe220786e4661b2bfda71ae41f7af388f03d;
mem[794] = 144'hf684fd3306a9e8aae19711271991115b1d9d;
mem[795] = 144'h1f39e553f8a3fd8fe6ba0d5d0501008a1c15;
mem[796] = 144'h1990edf0eab5e51c06edfe801893f4f812de;
mem[797] = 144'hf3970d841175103b04fe08c5eb61f478fa46;
mem[798] = 144'h0302e1cc0cdc0fe7f050187d155a09490364;
mem[799] = 144'hf4c0f4a10affeaf1175ef7300b35ef06045a;
mem[800] = 144'h08591357e7fa1150e91af1e1f74de744fa83;
mem[801] = 144'he69ffe78ff95161d02bdf46e11e00bb314dd;
mem[802] = 144'h17380480183de1d308bbf4461d84ff101e99;
mem[803] = 144'h126c0bb01f4b171c095114eb0cbdf9541e4e;
mem[804] = 144'h1e9e1593eae705a0f785183def13fd1fe319;
mem[805] = 144'he19f0eacf4b4fa4a094113e1e691ee681e4a;
mem[806] = 144'hf4dcea271c00ed7010650da4f0e2f7c61c77;
mem[807] = 144'h0a02099a0ac5151ef386f2a6ede7171de1e2;
mem[808] = 144'he521fa82fcb4f24cedfdff631e26e3c21390;
mem[809] = 144'hff7be92d17e61c5d0741f42ce97b09ba15d1;
mem[810] = 144'heb6e066e1dc60e85f5b9e5b3f14a11fa1477;
mem[811] = 144'hf639e5f7fc9809780dc1f398f988e7141fae;
mem[812] = 144'h00e304bbe34ee16116eaf9db097e11b6e36a;
mem[813] = 144'h109ef8b7e05afa96e9dc09b203db1b60e1b5;
mem[814] = 144'h1360e29be4321e7b00aaec40e5de1d35fc63;
mem[815] = 144'h1739e109ec83fa3515a4f257fe54e9d1f1a0;
mem[816] = 144'hea021ddb0be9f090fbad11151fc50c9d0e52;
mem[817] = 144'h017ffdaeea620790e1a8fda4fb900d8bfc26;
mem[818] = 144'hf12501fb190e1cabe30ff200e4d5e70de77e;
mem[819] = 144'hef74e3e8e867036300b81c8c021efa5d1aa3;
mem[820] = 144'h19e210c0e43a14a7e1b201befea018481a3e;
mem[821] = 144'hefec0db80de015c81571ff05f71efcca145e;
mem[822] = 144'h191c0553f4eb1816f506f2d0e5cf19bafd92;
mem[823] = 144'hea4df09de0a8ff0b16aa139610f31a2afb72;
mem[824] = 144'hf51ce5040104fcd1023e03f3e4ec0de2e35e;
mem[825] = 144'h0c06e0ebe609e0bdec21fddbf4b8ee4eefb4;
mem[826] = 144'h0bfcf557eb56e6501223f38c0d3ae2210a27;
mem[827] = 144'hf79a07cbe80eecf5e9e4f223e2baea34eab7;
mem[828] = 144'heeebf75f18451fb20062ed38e1a1052ce2b5;
mem[829] = 144'he3760d991c09ff33fafd05ba1103fa3f0044;
mem[830] = 144'h0397f468fbaae53d169819ef10340a46f04c;
mem[831] = 144'h0288ee0c1b631aa0031ef7a11ed1f9ca10d5;
mem[832] = 144'he0a6f18a006f07fce892e521f7e210301227;
mem[833] = 144'h08f0132afef5e59ee4a0f3ca137618afe7ea;
mem[834] = 144'h027a16f8edb31fc10cb2147d1bc41aa917a3;
mem[835] = 144'h0c8b0b4cfde8e1300a60085ced3411df09bb;
mem[836] = 144'he33e1f2ff8050ff10f54e82d1a16f643e7d0;
mem[837] = 144'h0da503a9ebca1aa5e308027fe08218cc16f6;
mem[838] = 144'hf7ad1d18e17ceee002a31c7c0b6dfa451c4c;
mem[839] = 144'h0cf80eae0f25f1981bf3ebd00ec30b460544;
mem[840] = 144'hf0710e8e0e1e12ba073ce7501174f31b191d;
mem[841] = 144'he230052b01591b7f11d5e8cee793e23eed5c;
mem[842] = 144'hec0bedcfe3a810acfa7ded1bfd8bf9d2e0f4;
mem[843] = 144'hf3f5e8d6f0061830011904d1e32b15b11aba;
mem[844] = 144'he04d182af50bfd320e83ee4cf88c03adeb8d;
mem[845] = 144'he7f4e943fd7b07e20485f4d3025cf0cfe175;
mem[846] = 144'hf982f814174c15be186fe455fe560bec1f3d;
mem[847] = 144'he4bc05791ac90b501c6f001ef0eb164a06e7;
mem[848] = 144'hf110e74bf61ce94ae6dff499f70aed6ff3d3;
mem[849] = 144'heab7f73d1939f131e7fc078de635fee81d4e;
mem[850] = 144'h034bfc91eaaf11e3f074f5e5f701fbb00458;
mem[851] = 144'he0faf3a7f7b10080eece00dcea0c19bbe712;
mem[852] = 144'hfa660d810e7d1b77f4cbed8a0a7bfbf3f6a2;
mem[853] = 144'h0ef0f85cfc2e051e05d9e0b3fdbde5ec1962;
mem[854] = 144'he0271639117afd5bfe9df9f81c411520f527;
mem[855] = 144'h04eff5b5f85efdbce43be1570b51f88be485;
mem[856] = 144'he4b616aa0e0214d61731e5cf11711fbd1016;
mem[857] = 144'he5d307ba0168f1aef404e606e601093d118d;
mem[858] = 144'h17a103f40cbe0d060f95e0c206f7ec89f8a7;
mem[859] = 144'h1fe11f0bffe715330192e8cff369125cf887;
mem[860] = 144'hf83ee7f10a0609d21a4def9718501069fe9a;
mem[861] = 144'hee721d90fded13af005fe344e3e00593f098;
mem[862] = 144'h0d4913691bad1da10b4ae4c9f245fd8cff4b;
mem[863] = 144'hffcb0333f301e21d1fdf07150702e4420147;
mem[864] = 144'h00c606861085f01af9d2024e0c11fb021886;
mem[865] = 144'h0a120f18e146edb709e41116f7d518f01e0d;
mem[866] = 144'h1da6f88d09691f520c3817e1e449fb5de7b1;
mem[867] = 144'h1130f64a0a160dac1ee30396f9be0ad600f0;
mem[868] = 144'hf3f2f612f8e701920a94eac5fbe3e866eed5;
mem[869] = 144'h19bbf6d1f75515de1f8606e1e790ffc5f32b;
mem[870] = 144'h10f4e585e56f19e7ede6e65ee9ce1e4d18e4;
mem[871] = 144'hf25fe9fd1ff00cfe0f10f898fe4617e80ba8;
mem[872] = 144'hf18bf60be39004f2e1e70343f45ae56b1aab;
mem[873] = 144'he02106da026ae606e561032a05a802e0f342;
mem[874] = 144'hf729185de7561830fb8f09b21a960630f94f;
mem[875] = 144'hea4ee560f137e6bffa83109f0f5ef92b1a94;
mem[876] = 144'h03cde591034e12391a2c115ef92ff333fefb;
mem[877] = 144'he25d1de7fa85e9ee16cb18791d5dec0eeab6;
mem[878] = 144'h0afb1d3e1393ee410a87fab5fb6908b10f66;
mem[879] = 144'hf44311c0010de45f0d6c0dd9ef3afd8ce602;
mem[880] = 144'h10890097ec2e04e2f7b51c1cf8e1f9f8156b;
mem[881] = 144'hec2a1c33e9fef429063a141ff1d60e1af177;
mem[882] = 144'hf141061aeb8bff34f73ef1271dd2e1e01e19;
mem[883] = 144'hf53e0e7f17e90ca8e5801f32fc01eaf8feca;
mem[884] = 144'hfb160268e24e0279ffddf6b416a809d103e3;
mem[885] = 144'h0256e559eda2f6d4f06aeeb30dfceea21852;
mem[886] = 144'hfb4f16e00248058912c9e2930ab503e8e209;
mem[887] = 144'he20af6f7ecf710d51357e829f03eeb5d17d2;
mem[888] = 144'h00a017e1f9af120d0433e611fa2be0f9e2bc;
mem[889] = 144'h1476f554ffe7144606fae89afe111fb411fd;
mem[890] = 144'h0e7afd67f0e916270bce0d2d09c209fee57d;
mem[891] = 144'h1f2504c3feabeab7e801e0bef3861481e23a;
mem[892] = 144'hfbfa1c7c1a38ff1d19b91794169df28f129b;
mem[893] = 144'hfc4b087de0d11fd1113d0b16e3b114e5151b;
mem[894] = 144'h099411ed1104e3ca1d1f0cacfb14e3be0116;
mem[895] = 144'hed3d1974e86d02ba0200e10803b7e1faf159;
mem[896] = 144'hf42c1cef140ee08af687fee5eba0eb9cfa28;
mem[897] = 144'he48c15541053f24cf25a0eeb15beee400b1c;
mem[898] = 144'hf0fff383e775e83102ae119f098f00aa15c2;
mem[899] = 144'hf4a1e6daf2df192dfa68081e1e67f477e45d;
mem[900] = 144'h1a8c0fa1e05d0ab516e4f755f959026604b1;
mem[901] = 144'hec1eed7e0223167ee6ca0c290ab9e716f055;
mem[902] = 144'he8551c551318e28c08d8f94912060bc40d94;
mem[903] = 144'hef95e0cae9951f72e4f8e18eed2ae6bee320;
mem[904] = 144'hf972149b1909f6c0e5d9e96a0359ecc500c4;
mem[905] = 144'h07381430035608c8f077f5801925face1947;
mem[906] = 144'h15f814fce0f4f4f919ed11e809eb00091fc9;
mem[907] = 144'he7b50968eda1ee1502d9e15ef6a3140f1039;
mem[908] = 144'h06ad061bfacf157e0d3ceb9a16201853f84c;
mem[909] = 144'h02cdf570ed5bf8fb1a6a1ca3fec20b5efb41;
mem[910] = 144'he4e30699f52a0077fd50e579fe3a1882e461;
mem[911] = 144'h0b98fecae6d0078a11ecfdf4f32ce5dde509;
mem[912] = 144'hfaa31ca51d0ee2f40f0dec371a82fb7d1188;
mem[913] = 144'h13101acf0472fc5ae77c192906ff0948f162;
mem[914] = 144'hf38de677f742fdb7ee3506c3fad61d97e3fb;
mem[915] = 144'h10f8f028f1760cd91ef5167d1b4ef15bf8e3;
mem[916] = 144'hf2381b7b09ff17c30fe9034ffdfe0eaaf361;
mem[917] = 144'h1082e54115421907ef7c00e203b9fccfec4c;
mem[918] = 144'h16821f71030bf1bf10d1064019ad02ee16cb;
mem[919] = 144'h09dfe03b13420e04fd54fa360387e934e482;
mem[920] = 144'he029ec300343e214f5b318d9fba1139e061d;
mem[921] = 144'hfb8af8ccec5104870cd2f56fe9791ca9ebf9;
mem[922] = 144'h16f906f0e561e674114915c31cccf051f9ba;
mem[923] = 144'hed92fec008a61e8fe614f59c03600ea3eb34;
mem[924] = 144'he588fa01fbc3f5be1d791783fa3e1c98f669;
mem[925] = 144'hef50f22d054502b5000fe754107df895ecaa;
mem[926] = 144'hea3c12e21bf91dc51478e72e05cff95ef03d;
mem[927] = 144'h099a1d440447f97ee0cce1a5e7ffe75be237;
mem[928] = 144'hefd5e2edeb1c1b25f37d08ad172a0784f9fa;
mem[929] = 144'hf36113a6042e1d0bfeb8dfcf1ccdf13a02fe;
mem[930] = 144'h03aef7c6f9bd0f8619f3e124062bf19af1cb;
mem[931] = 144'hf895fc17e52d1bfcff0dff5ff3b6eec51388;
mem[932] = 144'h04cce838102ceb9bf977e868fccde8751180;
mem[933] = 144'h078d105ffe3a0834f4a9ec83044ce209ebf1;
mem[934] = 144'hfe1413e01361f0160f58e0b400960ff1f281;
mem[935] = 144'heffbf8b11dccfd390bd4168e1167f4e5f7b3;
mem[936] = 144'he8250a33f99216d410fef0b1e77ffe0ce251;
mem[937] = 144'h1bfa184ffa6ce0031bb9ffffe4e01f5b1581;
mem[938] = 144'h1d280d22f8950c59fd790b251fa2eebbfb6b;
mem[939] = 144'h0a1d168d090d0ef71d0f16f4ec3a0296ec04;
mem[940] = 144'hfbba1f60101aff6e0b51f44fff4200cb0ddc;
mem[941] = 144'hfe260a0503ab04dfff86ea1cedaafc9e13bc;
mem[942] = 144'h0357ff83ebe6f56e003e162704551e2c06ed;
mem[943] = 144'he0690f74087efde5e565f08ef733f501ee3a;
mem[944] = 144'h0f63f8d7e94a0d4bf422019b1bfb1c33eae1;
mem[945] = 144'heba1fc3b17d9f8661a12f6f9096c0b15e907;
mem[946] = 144'hf834ee23e5b60b19f7e80ce0f62f0f89fa37;
mem[947] = 144'hedfe0594ebede0b20728e14317340cf51259;
mem[948] = 144'h139eee25e4540cbe00e70d77f4bc193be0e3;
mem[949] = 144'h1bb4e42d0874f98c03b515a9fdd0eef3171c;
mem[950] = 144'he0c8efdff432edc0e823f33af88d092d07b6;
mem[951] = 144'hfd9b18961af300e2e54beb3a04321428eba9;
mem[952] = 144'h1a97e55d1f19f5bd0395167310d7f3fae5f8;
mem[953] = 144'he17ce010ed24f31c0e340b00f4d1eca41793;
mem[954] = 144'h17d4e7ba18a0e56efc0c0bcf0996efe819fd;
mem[955] = 144'hf187f8a21fd2f1441971fa6c0585e1a4e918;
mem[956] = 144'h1d9d15edfbf7eef2012ae6bd1a9fe96ceae8;
mem[957] = 144'h029c1b42f8e8f9fbf71ff729fb94e1da0844;
mem[958] = 144'h136600eae322f4fa1e12f892f5f6096be119;
mem[959] = 144'h18740a74e9fbfd3f0c5b091e0567eee61dbc;
mem[960] = 144'hf54a1bb4f6bdfa60e2ecff3d07bb0b03fe82;
mem[961] = 144'h19ebf5581622e3eee5771b7ce6e71ce70c7f;
mem[962] = 144'hefba092a0bc217efe50be102edede779081d;
mem[963] = 144'h040df3a610a41476e0b7ef9a03daf3cee7ae;
mem[964] = 144'h0dfef4fef5b7ec17055cf6b817bcfd4ff119;
mem[965] = 144'hff6e0573ec99f010f2f7e63df7baff73fc74;
mem[966] = 144'h1c18f10bf9600b460bc7f63d101ee9561ebd;
mem[967] = 144'h14011c4e1136f6bb1c6be738006f0a40e40a;
mem[968] = 144'hf192091a11d2f954e965e26b0a59f2491e2a;
mem[969] = 144'heb9f1453eb7b184b02b1e124ed4d17ad0efa;
mem[970] = 144'hf9d1f3271bb900aae04b14220d19fb4a1dfe;
mem[971] = 144'hf4b9e40ff163f910ee230f02e2bbfb3a12ae;
mem[972] = 144'hef4f0a390c3df5321149f1a31a13e0dceb32;
mem[973] = 144'h1041f6141856f11b0b321f881b66fcd8ef06;
mem[974] = 144'he403f22d1becf2d3ff39f15ffa9cf635196d;
mem[975] = 144'heafc1412e2c91a7f133f01d8061f1510f2b9;
mem[976] = 144'h0b581fed0636135fec36f4e6f07eea7d0f10;
mem[977] = 144'he98de79e0c811a4ae5080064083105f81c7f;
mem[978] = 144'h0b4611b503011087e1fb0bc5e26c113d1ad3;
mem[979] = 144'hee1ffbdf1a37e2321130033502d41e54fa5e;
mem[980] = 144'h19acf5a4ffd5ecca0087096a1888e6711ba7;
mem[981] = 144'hf6cbf2201fd81fc30d5bf157e23ef608f8be;
mem[982] = 144'hf827e6c0fe1f036a0fd40c0bfd0415a2007c;
mem[983] = 144'hf3f1f533fbb8ff03e7cae8961be0ef2df4e8;
mem[984] = 144'h102003ff1ce01164188d021c17021ebdf42f;
mem[985] = 144'hfb61f6200a91fc1f198c0f62ed930caffa97;
mem[986] = 144'heeb60bb2ebe5fbfe16e2e038edfef3200ea2;
mem[987] = 144'hf9abebf5e38606f0e5abee331340123ce6bb;
mem[988] = 144'h0a65151ff0a1f76011f5f2fefae1e8cbf0eb;
mem[989] = 144'h0e20faff04a60821f240ec55e2b2167ee115;
mem[990] = 144'hf50efce102741a3f0dd5ff091dd2f30f03e5;
mem[991] = 144'h1d31f5ff19cdeaa9067de88beec51387fd9c;
mem[992] = 144'hef8412d4fa8913191424eb04e169ee72f850;
mem[993] = 144'h0f05fc8bf39a02ade54df0120532f31c099b;
mem[994] = 144'hf090fb681f1f0780081d182ce9b910f3fa92;
mem[995] = 144'hea68f3dc094101070f72e67c15e717321313;
mem[996] = 144'he38c1782f3f511570ef8fb38f5f4f9ab15a7;
mem[997] = 144'h13af0153e02608c9fbe2fc80174d05ce153f;
mem[998] = 144'h1781f28bf0e6ecfaf6eaf5820481e85413f1;
mem[999] = 144'heb35f897e3640d7a0d08e97afbaa0d181713;
mem[1000] = 144'h1e401a4d06c91c74e4560e581bae108604fd;
mem[1001] = 144'hedb0f3a406b2eea80f6d0e06e253ee6afe20;
mem[1002] = 144'hfde81028002bf211fb901840ec18e50a00ed;
mem[1003] = 144'h03f2f851f19205d30bef0b56f74100661286;
mem[1004] = 144'he985f1cbe51801bcf5da0dcd0b5bf6f31f2e;
mem[1005] = 144'h07f102b71ba70dabf798fa92f8ebf3f3f5bc;
mem[1006] = 144'h0f04181b1cfae5eee514109a12ab19001a8f;
mem[1007] = 144'he472f9d2eee90f78033e15551a341f450b8d;
mem[1008] = 144'h0c6ff76e026e16991eb1e056f7fd0a9bea24;
mem[1009] = 144'h1c7defa9e6b7f21bfcfbea0ce867f7bbec6c;
mem[1010] = 144'h1d8907bfed9ef1971bf8fba3f7e5029c0d89;
mem[1011] = 144'hf9941a9f011e09d0ede9fe5b126e07aaf02d;
mem[1012] = 144'h170c0b3f0b0201ea0ea110781d0d1792e177;
mem[1013] = 144'hf46b1e4707611048162804ba1d7ceedded37;
mem[1014] = 144'h17ddea5311c01f1cec33e81ef4b30bf10c1a;
mem[1015] = 144'h03d6ff2f1d71145d13ac0185106e110a0618;
mem[1016] = 144'h04b214e8ef81e80df535e06afe12e859ea5e;
mem[1017] = 144'h0c1cf2e9e2340ed2ff13efbc1ed806660906;
mem[1018] = 144'hfcd402e7e8920cac0d90fca2f237ecb8005f;
mem[1019] = 144'he72c0fe91c0cef8e09461a95efb00762eddc;
mem[1020] = 144'hf421e7c2f25e1cede7c5e66eea80e867e5b4;
mem[1021] = 144'hfc7d0bed0617f43cff7b1179f1071a1cf7a6;
mem[1022] = 144'h0e2eef15f8d8f32dfba1f7a31fad0536e163;
mem[1023] = 144'h0878f620fe0e047b0f93143e097a06d6ecbe;
mem[1024] = 144'hef1005e3ffb30ff1f8ac0c550e3c1806fcad;
mem[1025] = 144'h07b8e7d7142a019102fcec4a0e481d59f4d8;
mem[1026] = 144'hfff3f1e21ad6f587f47c086d1827eadd1e23;
mem[1027] = 144'he1500a240ce71046f973eb30025518490599;
mem[1028] = 144'he07fe11613bde04dec6def8df3d31d471dcd;
mem[1029] = 144'h1eaa0ba914be184feff3e6df1a3718f71976;
mem[1030] = 144'he1630f05ff9fe1d204c5021ef12e1c2ee258;
mem[1031] = 144'hee410779e9f90f3601650014fa920265fae8;
mem[1032] = 144'hfec3f6ea04970a3ee1bd122614c808270e07;
mem[1033] = 144'hf3d4f0071ef4ea8405011cc4edd3e132105d;
mem[1034] = 144'hfecb0e45f5b8047cf71414920951eb4d169e;
mem[1035] = 144'he85aed8c035af2c902e4138703ebfdb0f815;
mem[1036] = 144'he448f4161d51eb94041cf520e00319f116ec;
mem[1037] = 144'h0346f2a90288e8d10845fb9211c6f88413a6;
mem[1038] = 144'heee10024133ff8a40e8c038de185e9d710bb;
mem[1039] = 144'h04f2034ffca5f404190efc9ee368133e0490;
mem[1040] = 144'h0711f9bafb61174a0eedfb630efa17ce07ff;
mem[1041] = 144'h037210e2e4cb1dcaead2ec1dfebf03b0f5e9;
mem[1042] = 144'hfb35fe950a8f157c0faf057ffc361b83fbde;
mem[1043] = 144'hfb15eb52e2e2f1e9f0cbf4d0e01df3a7e25a;
mem[1044] = 144'h0df2011e0b521d24fd1dec0f1b9ee15ff977;
mem[1045] = 144'hf84ef9b5fa7ffda5148be72a10740451fd68;
mem[1046] = 144'h17edfc55081f09a3f0c819de0ec6fd24e736;
mem[1047] = 144'hec76e72ae8fe1ca803b4040d11bdea050021;
mem[1048] = 144'he79010e10dd0e4e0f1edfa74e5b2fd42e189;
mem[1049] = 144'hfcc21489ef8c042f1939e74df9b00da31a16;
mem[1050] = 144'heb4bfd950553002f11fb15080756e53afa54;
mem[1051] = 144'he4b3fc65030f1450f0f6073b08030704e773;
mem[1052] = 144'hefd5f6e716a4ea1aee0f175205de1e72f8c0;
mem[1053] = 144'hed79f5b7f475f322fefa0acd1e87fa8b01e0;
mem[1054] = 144'h03f50525e3f9fd27f603e6aee339e0cb10f6;
mem[1055] = 144'he044e7171f47e473e6aa15fd1dbb0ed4e385;
mem[1056] = 144'hffb60043edc2f4f2186c1cd3eba41a700edd;
mem[1057] = 144'hf4ee0163f2bb0ccfe419f5e9fd21fec313d9;
mem[1058] = 144'h045af41b0f96f8b2f27eee9208d3ed5408aa;
mem[1059] = 144'he036094918fa0699e509e711f7b108140ba0;
mem[1060] = 144'h0d7f00c91b9118250131e9c6ea5d1c7a00fa;
mem[1061] = 144'he5c6e6531954f19214d9e109f24c1524ea76;
mem[1062] = 144'h17b30f7500c9e639f913f218e077e7211f2a;
mem[1063] = 144'hf3c1f3a70dc4f6741afdfc63f9f9ef22f66a;
mem[1064] = 144'h03140ef90388fb93ed3eec28f3240b48f5ee;
mem[1065] = 144'he915f00bf0f009efe2d9e8a7e3c30145f196;
mem[1066] = 144'hf843e2b7ed98e34706c217d917cb08fe0493;
mem[1067] = 144'heb58ec9c105a1c22e02c03d1f3550c05e054;
mem[1068] = 144'hfb97eb26e1ae01e7f637018a1309ed20f12a;
mem[1069] = 144'he442f11f1f9ff82700951eaf18a30aadebc8;
mem[1070] = 144'h13fff36ef377e6df0d791ed7ff2b1db1f275;
mem[1071] = 144'hfd5b14c9eea518b5e533e5dc1d5711540a0f;
mem[1072] = 144'hf2a8f2fff843f97ee0df1668e6500a51ec46;
mem[1073] = 144'hfadfeef813a61c9aeea8f309fbdd13df15b5;
mem[1074] = 144'h073c14f0f839e524e7f51238f8d2e14419b3;
mem[1075] = 144'he2dfe2420b0c18e2ee16fb68fbe9089314eb;
mem[1076] = 144'heb3cf95908e417d4e98b1f701cfd1b010ed3;
mem[1077] = 144'he159fa8d00c5fe57f053fb3af51deabef133;
mem[1078] = 144'he6dc1ff2160cf87ff48c01c4097ee3f1f09e;
mem[1079] = 144'h09c712e41c850abe1dabfac7f678ec5ae83f;
mem[1080] = 144'h0ccae524f8e61c4f115a0acfe5120d43ff04;
mem[1081] = 144'h13f6f9e61276e29fe82be996fc990eccf761;
mem[1082] = 144'hf780e33bf7421a6c02aff19bf1e7ee8cf02d;
mem[1083] = 144'hec00f28d064de4cc0526f7ddfe3fefdb1ac7;
mem[1084] = 144'h0cde1c72fcb91d1fe0cbf7c01608e5221258;
mem[1085] = 144'he84911b318670d0d0da2e717e702f2760923;
mem[1086] = 144'he756e87f0c6108b5fec7101c126600e50079;
mem[1087] = 144'h0cbaead2e8d411870e99fba415fe01bbe350;
mem[1088] = 144'hef97eae21696efa70e95e68eeac1eac2f7f4;
mem[1089] = 144'hfe11fee6f678ef89e5bc1b69e3db15a118d6;
mem[1090] = {16'h0978, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1091] = {16'h0434, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1092] = {16'h03d5, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1093] = {16'h11fd, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1094] = {16'he72f, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1095] = {16'heb72, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1096] = {16'hf186, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1097] = {16'h0e24, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1098] = {16'h1738, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
mem[1099] = {16'h02b9, 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule