// Module: top.sv
// Date: 11/1/2019
// Description: Top level module. Wraps the controller (core of the CNN) and RAM elements.

`timescale 1ns/1ns

module top #(parameter 
    GS_BITS = 8, 
    BCD_BITS = 4, 
    D_WIDTH = 16,

    LINE_BUF_GROUPS = 16,
    LINE_BUFS_PER_GROUP = 2,
    LINE_BUF_DEPTH = 30,
    LINE_BUF_ADDR_BITS = 5,
    
    FMAP_I_MEM_BLKS = 16,
    FMAP_I_DEPTH = 196,
    FMAP_I_ADDR_BITS = 8,

    FMAP_II_MEM_BLKS = 144,
    FMAP_II_DEPTH = 8,
    FMAP_II_ADDR_BITS = 3,

    FMAP_III_MEM_BLKS = 64,
    FMAP_III_DEPTH = 1,
    FMAP_III_ADDR_BITS = 1,

    WEIGHT_MEM_BLKS = 16,
    WEIGHT_MEM_DEPTH = 1100,
    WEIGHT_MEM_ADDR_BITS = 11,
    WEIGHT_MEM_D_WIDTH = 144,

    BIAS_MEM_DEPTH = 16,
    BIAS_MEM_ADDR_BITS = 4,
    BIAS_MEM_D_WIDTH = 128

) (
    // input MNIST image to the convolutional neural network
    input clk,
    input rst,
    input [GS_BITS-1:0] pixel_i,
    input pixel_i_valid, 

    // digit classification output
    output reg [BCD_BITS-1:0] digit_o,
    output reg digit_o_valid
    
);

// Line buffers
wire [D_WIDTH-1:0] line_buffer_rd_data [LINE_BUF_GROUPS-1:0][LINE_BUFS_PER_GROUP-1:0]; // 16-b data
wire [LINE_BUF_ADDR_BITS-1:0] line_buffer_rd_addr [LINE_BUF_GROUPS-1:0][LINE_BUFS_PER_GROUP-1:0]; // log2(30) = 5 bits
wire [LINE_BUF_ADDR_BITS-1:0] line_buffer_wr_addr [LINE_BUF_GROUPS-1:0][LINE_BUFS_PER_GROUP-1:0];
wire [D_WIDTH-1:0] line_buffer_wr_data [LINE_BUF_GROUPS-1:0][LINE_BUFS_PER_GROUP-1:0];
wire line_buffer_wr_en [LINE_BUF_GROUPS-1:0][LINE_BUFS_PER_GROUP-1:0];

// fmap I memory I/O, for the resulting fmaps of CONV2. (input image -> CONV2 -> fmap I)
wire [FMAP_I_ADDR_BITS-1:0] fmap_wr_addr_I [FMAP_I_MEM_BLKS-1:0]; 
wire [FMAP_I_ADDR_BITS-1:0] fmap_rd_addr_I [FMAP_I_MEM_BLKS-1:0];
wire fmap_wr_en_I [FMAP_I_MEM_BLKS-1:0];
wire [D_WIDTH-1:0] fmap_wr_data_I [FMAP_I_MEM_BLKS-1:0];
wire [D_WIDTH-1:0] fmap_rd_data_I [FMAP_I_MEM_BLKS-1:0];

// fmap II memory I/O, for the resulting fmaps of CONV4. (fmap I -> CONV4 -> fmap II)
wire [FMAP_II_ADDR_BITS-1:0] fmap_wr_addr_II [FMAP_II_MEM_BLKS-1:0];
wire [FMAP_II_ADDR_BITS-1:0] fmap_rd_addr_II [FMAP_II_MEM_BLKS-1:0];
wire fmap_wr_en_II [FMAP_II_MEM_BLKS-1:0];
wire [D_WIDTH-1:0] fmap_wr_data_II [FMAP_II_MEM_BLKS-1:0];
wire [D_WIDTH-1:0] fmap_rd_data_II [FMAP_II_MEM_BLKS-1:0];

// fmap III memory I/O, for the resulting fmaps of FC6. (fmap II -> FC6 -> fmap III).
wire [FMAP_III_ADDR_BITS-1:0] fmap_wr_addr_III [FMAP_III_MEM_BLKS-1:0];
wire [FMAP_III_ADDR_BITS-1:0] fmap_rd_addr_III [FMAP_III_MEM_BLKS-1:0];
wire fmap_wr_en_III [FMAP_III_MEM_BLKS-1:0];
wire [D_WIDTH-1:0] fmap_wr_data_III [FMAP_III_MEM_BLKS-1:0];
wire [D_WIDTH-1:0] fmap_rd_data_III [FMAP_III_MEM_BLKS-1:0];

// Weight memory (dual port ROM)
wire [WEIGHT_MEM_ADDR_BITS-1:0] addr_a [WEIGHT_MEM_BLKS/2-1:0];
wire [WEIGHT_MEM_ADDR_BITS-1:0] addr_b [WEIGHT_MEM_BLKS/2-1:0];
wire [WEIGHT_MEM_D_WIDTH-1:0] q_a [WEIGHT_MEM_BLKS/2-1:0];
wire [WEIGHT_MEM_D_WIDTH-1:0] q_b [WEIGHT_MEM_BLKS/2-1:0];

// Bias memory (dual port ROM)
wire [BIAS_MEM_ADDR_BITS-1:0] bi_addr_a;
wire [BIAS_MEM_ADDR_BITS-1:0] bi_addr_b;
wire [BIAS_MEM_D_WIDTH-1:0] bi_q_a;
wire [BIAS_MEM_D_WIDTH-1:0] bi_q_b;

// CNN core
controller controller_u 
(
    .clk       (clk),
    .rst       (rst),

    // Ifmap pixel input
    .pixel_i       (pixel_i),
    .pixel_i_valid (pixel_i_valid),

    // Weights I/O
    .\addr_a[0]  (addr_a[0] ),
    .\addr_a[1]  (addr_a[1] ),
    .\addr_a[2]  (addr_a[2] ),
    .\addr_a[3]  (addr_a[3] ),
    .\addr_a[4]  (addr_a[4] ),
    .\addr_a[5]  (addr_a[5] ),
    .\addr_a[6]  (addr_a[6] ),
    .\addr_a[7]  (addr_a[7] ),

    .\addr_b[0]  (addr_b[0] ),
    .\addr_b[1]  (addr_b[1] ),
    .\addr_b[2]  (addr_b[2] ),
    .\addr_b[3]  (addr_b[3] ),
    .\addr_b[4]  (addr_b[4] ),
    .\addr_b[5]  (addr_b[5] ),
    .\addr_b[6]  (addr_b[6] ),
    .\addr_b[7]  (addr_b[7] ),

    .\q_a[0]  (q_a[0] ),
    .\q_a[1]  (q_a[1] ),
    .\q_a[2]  (q_a[2] ),
    .\q_a[3]  (q_a[3] ),
    .\q_a[4]  (q_a[4] ),
    .\q_a[5]  (q_a[5] ),
    .\q_a[6]  (q_a[6] ),
    .\q_a[7]  (q_a[7] ),

    .\q_b[0]  (q_b[0] ),
    .\q_b[1]  (q_b[1] ),
    .\q_b[2]  (q_b[2] ),
    .\q_b[3]  (q_b[3] ),
    .\q_b[4]  (q_b[4] ),
    .\q_b[5]  (q_b[5] ),
    .\q_b[6]  (q_b[6] ),
    .\q_b[7]  (q_b[7] ),

    .bi_addr_a  (bi_addr_a),
    .bi_addr_b  (bi_addr_b),
    .bi_q_a     (bi_q_a),
    .bi_q_b     (bi_q_b),

    .\line_buffer_rd_data[0][0]	(line_buffer_rd_data[0][0]	),
    .\line_buffer_rd_data[0][1]	(line_buffer_rd_data[0][1]	),
    .\line_buffer_rd_data[1][0]	(line_buffer_rd_data[1][0]	),
    .\line_buffer_rd_data[1][1]	(line_buffer_rd_data[1][1]	),
    .\line_buffer_rd_data[2][0]	(line_buffer_rd_data[2][0]	),
    .\line_buffer_rd_data[2][1]	(line_buffer_rd_data[2][1]	),
    .\line_buffer_rd_data[3][0]	(line_buffer_rd_data[3][0]	),
    .\line_buffer_rd_data[3][1]	(line_buffer_rd_data[3][1]	),
    .\line_buffer_rd_data[4][0]	(line_buffer_rd_data[4][0]	),
    .\line_buffer_rd_data[4][1]	(line_buffer_rd_data[4][1]	),
    .\line_buffer_rd_data[5][0]	(line_buffer_rd_data[5][0]	),
    .\line_buffer_rd_data[5][1]	(line_buffer_rd_data[5][1]	),
    .\line_buffer_rd_data[6][0]	(line_buffer_rd_data[6][0]	),
    .\line_buffer_rd_data[6][1]	(line_buffer_rd_data[6][1]	),
    .\line_buffer_rd_data[7][0]	(line_buffer_rd_data[7][0]	),
    .\line_buffer_rd_data[7][1]	(line_buffer_rd_data[7][1]	),
    .\line_buffer_rd_data[8][0]	(line_buffer_rd_data[8][0]	),
    .\line_buffer_rd_data[8][1]	(line_buffer_rd_data[8][1]	),
    .\line_buffer_rd_data[9][0]	(line_buffer_rd_data[9][0]	),
    .\line_buffer_rd_data[9][1]	(line_buffer_rd_data[9][1]	),
    .\line_buffer_rd_data[10][0]	(line_buffer_rd_data[10][0]	),
    .\line_buffer_rd_data[10][1]	(line_buffer_rd_data[10][1]	),
    .\line_buffer_rd_data[11][0]	(line_buffer_rd_data[11][0]	),
    .\line_buffer_rd_data[11][1]	(line_buffer_rd_data[11][1]	),
    .\line_buffer_rd_data[12][0]	(line_buffer_rd_data[12][0]	),
    .\line_buffer_rd_data[12][1]	(line_buffer_rd_data[12][1]	),
    .\line_buffer_rd_data[13][0]	(line_buffer_rd_data[13][0]	),
    .\line_buffer_rd_data[13][1]	(line_buffer_rd_data[13][1]	),
    .\line_buffer_rd_data[14][0]	(line_buffer_rd_data[14][0]	),
    .\line_buffer_rd_data[14][1]	(line_buffer_rd_data[14][1]	),
    .\line_buffer_rd_data[15][0]	(line_buffer_rd_data[15][0]	),
    .\line_buffer_rd_data[15][1]	(line_buffer_rd_data[15][1]	),

    .\line_buffer_rd_addr[0][0]	(line_buffer_rd_addr[0][0]	),
    .\line_buffer_rd_addr[0][1]	(line_buffer_rd_addr[0][1]	),
    .\line_buffer_rd_addr[1][0]	(line_buffer_rd_addr[1][0]	),
    .\line_buffer_rd_addr[1][1]	(line_buffer_rd_addr[1][1]	),
    .\line_buffer_rd_addr[2][0]	(line_buffer_rd_addr[2][0]	),
    .\line_buffer_rd_addr[2][1]	(line_buffer_rd_addr[2][1]	),
    .\line_buffer_rd_addr[3][0]	(line_buffer_rd_addr[3][0]	),
    .\line_buffer_rd_addr[3][1]	(line_buffer_rd_addr[3][1]	),
    .\line_buffer_rd_addr[4][0]	(line_buffer_rd_addr[4][0]	),
    .\line_buffer_rd_addr[4][1]	(line_buffer_rd_addr[4][1]	),
    .\line_buffer_rd_addr[5][0]	(line_buffer_rd_addr[5][0]	),
    .\line_buffer_rd_addr[5][1]	(line_buffer_rd_addr[5][1]	),
    .\line_buffer_rd_addr[6][0]	(line_buffer_rd_addr[6][0]	),
    .\line_buffer_rd_addr[6][1]	(line_buffer_rd_addr[6][1]	),
    .\line_buffer_rd_addr[7][0]	(line_buffer_rd_addr[7][0]	),
    .\line_buffer_rd_addr[7][1]	(line_buffer_rd_addr[7][1]	),
    .\line_buffer_rd_addr[8][0]	(line_buffer_rd_addr[8][0]	),
    .\line_buffer_rd_addr[8][1]	(line_buffer_rd_addr[8][1]	),
    .\line_buffer_rd_addr[9][0]	(line_buffer_rd_addr[9][0]	),
    .\line_buffer_rd_addr[9][1]	(line_buffer_rd_addr[9][1]	),
    .\line_buffer_rd_addr[10][0]	(line_buffer_rd_addr[10][0]	),
    .\line_buffer_rd_addr[10][1]	(line_buffer_rd_addr[10][1]	),
    .\line_buffer_rd_addr[11][0]	(line_buffer_rd_addr[11][0]	),
    .\line_buffer_rd_addr[11][1]	(line_buffer_rd_addr[11][1]	),
    .\line_buffer_rd_addr[12][0]	(line_buffer_rd_addr[12][0]	),
    .\line_buffer_rd_addr[12][1]	(line_buffer_rd_addr[12][1]	),
    .\line_buffer_rd_addr[13][0]	(line_buffer_rd_addr[13][0]	),
    .\line_buffer_rd_addr[13][1]	(line_buffer_rd_addr[13][1]	),
    .\line_buffer_rd_addr[14][0]	(line_buffer_rd_addr[14][0]	),
    .\line_buffer_rd_addr[14][1]	(line_buffer_rd_addr[14][1]	),
    .\line_buffer_rd_addr[15][0]	(line_buffer_rd_addr[15][0]	),
    .\line_buffer_rd_addr[15][1]	(line_buffer_rd_addr[15][1]	),

    .\line_buffer_wr_addr[0][0]	(line_buffer_wr_addr[0][0]	),
    .\line_buffer_wr_addr[0][1]	(line_buffer_wr_addr[0][1]	),
    .\line_buffer_wr_addr[1][0]	(line_buffer_wr_addr[1][0]	),
    .\line_buffer_wr_addr[1][1]	(line_buffer_wr_addr[1][1]	),
    .\line_buffer_wr_addr[2][0]	(line_buffer_wr_addr[2][0]	),
    .\line_buffer_wr_addr[2][1]	(line_buffer_wr_addr[2][1]	),
    .\line_buffer_wr_addr[3][0]	(line_buffer_wr_addr[3][0]	),
    .\line_buffer_wr_addr[3][1]	(line_buffer_wr_addr[3][1]	),
    .\line_buffer_wr_addr[4][0]	(line_buffer_wr_addr[4][0]	),
    .\line_buffer_wr_addr[4][1]	(line_buffer_wr_addr[4][1]	),
    .\line_buffer_wr_addr[5][0]	(line_buffer_wr_addr[5][0]	),
    .\line_buffer_wr_addr[5][1]	(line_buffer_wr_addr[5][1]	),
    .\line_buffer_wr_addr[6][0]	(line_buffer_wr_addr[6][0]	),
    .\line_buffer_wr_addr[6][1]	(line_buffer_wr_addr[6][1]	),
    .\line_buffer_wr_addr[7][0]	(line_buffer_wr_addr[7][0]	),
    .\line_buffer_wr_addr[7][1]	(line_buffer_wr_addr[7][1]	),
    .\line_buffer_wr_addr[8][0]	(line_buffer_wr_addr[8][0]	),
    .\line_buffer_wr_addr[8][1]	(line_buffer_wr_addr[8][1]	),
    .\line_buffer_wr_addr[9][0]	(line_buffer_wr_addr[9][0]	),
    .\line_buffer_wr_addr[9][1]	(line_buffer_wr_addr[9][1]	),
    .\line_buffer_wr_addr[10][0]	(line_buffer_wr_addr[10][0]	),
    .\line_buffer_wr_addr[10][1]	(line_buffer_wr_addr[10][1]	),
    .\line_buffer_wr_addr[11][0]	(line_buffer_wr_addr[11][0]	),
    .\line_buffer_wr_addr[11][1]	(line_buffer_wr_addr[11][1]	),
    .\line_buffer_wr_addr[12][0]	(line_buffer_wr_addr[12][0]	),
    .\line_buffer_wr_addr[12][1]	(line_buffer_wr_addr[12][1]	),
    .\line_buffer_wr_addr[13][0]	(line_buffer_wr_addr[13][0]	),
    .\line_buffer_wr_addr[13][1]	(line_buffer_wr_addr[13][1]	),
    .\line_buffer_wr_addr[14][0]	(line_buffer_wr_addr[14][0]	),
    .\line_buffer_wr_addr[14][1]	(line_buffer_wr_addr[14][1]	),
    .\line_buffer_wr_addr[15][0]	(line_buffer_wr_addr[15][0]	),
    .\line_buffer_wr_addr[15][1]	(line_buffer_wr_addr[15][1]	),

    .\line_buffer_wr_data[0][0]	(line_buffer_wr_data[0][0]	),
    .\line_buffer_wr_data[0][1]	(line_buffer_wr_data[0][1]	),
    .\line_buffer_wr_data[1][0]	(line_buffer_wr_data[1][0]	),
    .\line_buffer_wr_data[1][1]	(line_buffer_wr_data[1][1]	),
    .\line_buffer_wr_data[2][0]	(line_buffer_wr_data[2][0]	),
    .\line_buffer_wr_data[2][1]	(line_buffer_wr_data[2][1]	),
    .\line_buffer_wr_data[3][0]	(line_buffer_wr_data[3][0]	),
    .\line_buffer_wr_data[3][1]	(line_buffer_wr_data[3][1]	),
    .\line_buffer_wr_data[4][0]	(line_buffer_wr_data[4][0]	),
    .\line_buffer_wr_data[4][1]	(line_buffer_wr_data[4][1]	),
    .\line_buffer_wr_data[5][0]	(line_buffer_wr_data[5][0]	),
    .\line_buffer_wr_data[5][1]	(line_buffer_wr_data[5][1]	),
    .\line_buffer_wr_data[6][0]	(line_buffer_wr_data[6][0]	),
    .\line_buffer_wr_data[6][1]	(line_buffer_wr_data[6][1]	),
    .\line_buffer_wr_data[7][0]	(line_buffer_wr_data[7][0]	),
    .\line_buffer_wr_data[7][1]	(line_buffer_wr_data[7][1]	),
    .\line_buffer_wr_data[8][0]	(line_buffer_wr_data[8][0]	),
    .\line_buffer_wr_data[8][1]	(line_buffer_wr_data[8][1]	),
    .\line_buffer_wr_data[9][0]	(line_buffer_wr_data[9][0]	),
    .\line_buffer_wr_data[9][1]	(line_buffer_wr_data[9][1]	),
    .\line_buffer_wr_data[10][0]	(line_buffer_wr_data[10][0]	),
    .\line_buffer_wr_data[10][1]	(line_buffer_wr_data[10][1]	),
    .\line_buffer_wr_data[11][0]	(line_buffer_wr_data[11][0]	),
    .\line_buffer_wr_data[11][1]	(line_buffer_wr_data[11][1]	),
    .\line_buffer_wr_data[12][0]	(line_buffer_wr_data[12][0]	),
    .\line_buffer_wr_data[12][1]	(line_buffer_wr_data[12][1]	),
    .\line_buffer_wr_data[13][0]	(line_buffer_wr_data[13][0]	),
    .\line_buffer_wr_data[13][1]	(line_buffer_wr_data[13][1]	),
    .\line_buffer_wr_data[14][0]	(line_buffer_wr_data[14][0]	),
    .\line_buffer_wr_data[14][1]	(line_buffer_wr_data[14][1]	),
    .\line_buffer_wr_data[15][0]	(line_buffer_wr_data[15][0]	),
    .\line_buffer_wr_data[15][1]	(line_buffer_wr_data[15][1]	),

    .\line_buffer_wr_en[0][0]	(line_buffer_wr_en[0][0]	),
    .\line_buffer_wr_en[0][1]	(line_buffer_wr_en[0][1]	),
    .\line_buffer_wr_en[1][0]	(line_buffer_wr_en[1][0]	),
    .\line_buffer_wr_en[1][1]	(line_buffer_wr_en[1][1]	),
    .\line_buffer_wr_en[2][0]	(line_buffer_wr_en[2][0]	),
    .\line_buffer_wr_en[2][1]	(line_buffer_wr_en[2][1]	),
    .\line_buffer_wr_en[3][0]	(line_buffer_wr_en[3][0]	),
    .\line_buffer_wr_en[3][1]	(line_buffer_wr_en[3][1]	),
    .\line_buffer_wr_en[4][0]	(line_buffer_wr_en[4][0]	),
    .\line_buffer_wr_en[4][1]	(line_buffer_wr_en[4][1]	),
    .\line_buffer_wr_en[5][0]	(line_buffer_wr_en[5][0]	),
    .\line_buffer_wr_en[5][1]	(line_buffer_wr_en[5][1]	),
    .\line_buffer_wr_en[6][0]	(line_buffer_wr_en[6][0]	),
    .\line_buffer_wr_en[6][1]	(line_buffer_wr_en[6][1]	),
    .\line_buffer_wr_en[7][0]	(line_buffer_wr_en[7][0]	),
    .\line_buffer_wr_en[7][1]	(line_buffer_wr_en[7][1]	),
    .\line_buffer_wr_en[8][0]	(line_buffer_wr_en[8][0]	),
    .\line_buffer_wr_en[8][1]	(line_buffer_wr_en[8][1]	),
    .\line_buffer_wr_en[9][0]	(line_buffer_wr_en[9][0]	),
    .\line_buffer_wr_en[9][1]	(line_buffer_wr_en[9][1]	),
    .\line_buffer_wr_en[10][0]	(line_buffer_wr_en[10][0]	),
    .\line_buffer_wr_en[10][1]	(line_buffer_wr_en[10][1]	),
    .\line_buffer_wr_en[11][0]	(line_buffer_wr_en[11][0]	),
    .\line_buffer_wr_en[11][1]	(line_buffer_wr_en[11][1]	),
    .\line_buffer_wr_en[12][0]	(line_buffer_wr_en[12][0]	),
    .\line_buffer_wr_en[12][1]	(line_buffer_wr_en[12][1]	),
    .\line_buffer_wr_en[13][0]	(line_buffer_wr_en[13][0]	),
    .\line_buffer_wr_en[13][1]	(line_buffer_wr_en[13][1]	),
    .\line_buffer_wr_en[14][0]	(line_buffer_wr_en[14][0]	),
    .\line_buffer_wr_en[14][1]	(line_buffer_wr_en[14][1]	),
    .\line_buffer_wr_en[15][0]	(line_buffer_wr_en[15][0]	),
    .\line_buffer_wr_en[15][1]	(line_buffer_wr_en[15][1]	),

    .\fmap_wr_addr_I[0]	(fmap_wr_addr_I[0]	),
    .\fmap_wr_addr_I[1]	(fmap_wr_addr_I[1]	),
    .\fmap_wr_addr_I[2]	(fmap_wr_addr_I[2]	),
    .\fmap_wr_addr_I[3]	(fmap_wr_addr_I[3]	),
    .\fmap_wr_addr_I[4]	(fmap_wr_addr_I[4]	),
    .\fmap_wr_addr_I[5]	(fmap_wr_addr_I[5]	),
    .\fmap_wr_addr_I[6]	(fmap_wr_addr_I[6]	),
    .\fmap_wr_addr_I[7]	(fmap_wr_addr_I[7]	),
    .\fmap_wr_addr_I[8]	(fmap_wr_addr_I[8]	),
    .\fmap_wr_addr_I[9]	(fmap_wr_addr_I[9]	),
    .\fmap_wr_addr_I[10]	(fmap_wr_addr_I[10]	),
    .\fmap_wr_addr_I[11]	(fmap_wr_addr_I[11]	),
    .\fmap_wr_addr_I[12]	(fmap_wr_addr_I[12]	),
    .\fmap_wr_addr_I[13]	(fmap_wr_addr_I[13]	),
    .\fmap_wr_addr_I[14]	(fmap_wr_addr_I[14]	),
    .\fmap_wr_addr_I[15]	(fmap_wr_addr_I[15]	),

    .\fmap_rd_addr_I[0]	(fmap_rd_addr_I[0]	),
    .\fmap_rd_addr_I[1]	(fmap_rd_addr_I[1]	),
    .\fmap_rd_addr_I[2]	(fmap_rd_addr_I[2]	),
    .\fmap_rd_addr_I[3]	(fmap_rd_addr_I[3]	),
    .\fmap_rd_addr_I[4]	(fmap_rd_addr_I[4]	),
    .\fmap_rd_addr_I[5]	(fmap_rd_addr_I[5]	),
    .\fmap_rd_addr_I[6]	(fmap_rd_addr_I[6]	),
    .\fmap_rd_addr_I[7]	(fmap_rd_addr_I[7]	),
    .\fmap_rd_addr_I[8]	(fmap_rd_addr_I[8]	),
    .\fmap_rd_addr_I[9]	(fmap_rd_addr_I[9]	),
    .\fmap_rd_addr_I[10]	(fmap_rd_addr_I[10]	),
    .\fmap_rd_addr_I[11]	(fmap_rd_addr_I[11]	),
    .\fmap_rd_addr_I[12]	(fmap_rd_addr_I[12]	),
    .\fmap_rd_addr_I[13]	(fmap_rd_addr_I[13]	),
    .\fmap_rd_addr_I[14]	(fmap_rd_addr_I[14]	),
    .\fmap_rd_addr_I[15]	(fmap_rd_addr_I[15]	),

    .\fmap_wr_en_I[0]	(fmap_wr_en_I[0]	),
    .\fmap_wr_en_I[1]	(fmap_wr_en_I[1]	),
    .\fmap_wr_en_I[2]	(fmap_wr_en_I[2]	),
    .\fmap_wr_en_I[3]	(fmap_wr_en_I[3]	),
    .\fmap_wr_en_I[4]	(fmap_wr_en_I[4]	),
    .\fmap_wr_en_I[5]	(fmap_wr_en_I[5]	),
    .\fmap_wr_en_I[6]	(fmap_wr_en_I[6]	),
    .\fmap_wr_en_I[7]	(fmap_wr_en_I[7]	),
    .\fmap_wr_en_I[8]	(fmap_wr_en_I[8]	),
    .\fmap_wr_en_I[9]	(fmap_wr_en_I[9]	),
    .\fmap_wr_en_I[10]	(fmap_wr_en_I[10]	),
    .\fmap_wr_en_I[11]	(fmap_wr_en_I[11]	),
    .\fmap_wr_en_I[12]	(fmap_wr_en_I[12]	),
    .\fmap_wr_en_I[13]	(fmap_wr_en_I[13]	),
    .\fmap_wr_en_I[14]	(fmap_wr_en_I[14]	),
    .\fmap_wr_en_I[15]	(fmap_wr_en_I[15]	),

    .\fmap_wr_data_I[0]	(fmap_wr_data_I[0]	),
    .\fmap_wr_data_I[1]	(fmap_wr_data_I[1]	),
    .\fmap_wr_data_I[2]	(fmap_wr_data_I[2]	),
    .\fmap_wr_data_I[3]	(fmap_wr_data_I[3]	),
    .\fmap_wr_data_I[4]	(fmap_wr_data_I[4]	),
    .\fmap_wr_data_I[5]	(fmap_wr_data_I[5]	),
    .\fmap_wr_data_I[6]	(fmap_wr_data_I[6]	),
    .\fmap_wr_data_I[7]	(fmap_wr_data_I[7]	),
    .\fmap_wr_data_I[8]	(fmap_wr_data_I[8]	),
    .\fmap_wr_data_I[9]	(fmap_wr_data_I[9]	),
    .\fmap_wr_data_I[10]	(fmap_wr_data_I[10]	),
    .\fmap_wr_data_I[11]	(fmap_wr_data_I[11]	),
    .\fmap_wr_data_I[12]	(fmap_wr_data_I[12]	),
    .\fmap_wr_data_I[13]	(fmap_wr_data_I[13]	),
    .\fmap_wr_data_I[14]	(fmap_wr_data_I[14]	),
    .\fmap_wr_data_I[15]	(fmap_wr_data_I[15]	),

    .\fmap_rd_data_I[0]	(fmap_rd_data_I[0]	),
    .\fmap_rd_data_I[1]	(fmap_rd_data_I[1]	),
    .\fmap_rd_data_I[2]	(fmap_rd_data_I[2]	),
    .\fmap_rd_data_I[3]	(fmap_rd_data_I[3]	),
    .\fmap_rd_data_I[4]	(fmap_rd_data_I[4]	),
    .\fmap_rd_data_I[5]	(fmap_rd_data_I[5]	),
    .\fmap_rd_data_I[6]	(fmap_rd_data_I[6]	),
    .\fmap_rd_data_I[7]	(fmap_rd_data_I[7]	),
    .\fmap_rd_data_I[8]	(fmap_rd_data_I[8]	),
    .\fmap_rd_data_I[9]	(fmap_rd_data_I[9]	),
    .\fmap_rd_data_I[10]	(fmap_rd_data_I[10]	),
    .\fmap_rd_data_I[11]	(fmap_rd_data_I[11]	),
    .\fmap_rd_data_I[12]	(fmap_rd_data_I[12]	),
    .\fmap_rd_data_I[13]	(fmap_rd_data_I[13]	),
    .\fmap_rd_data_I[14]	(fmap_rd_data_I[14]	),
    .\fmap_rd_data_I[15]	(fmap_rd_data_I[15]	),

    .\fmap_rd_data_II[0]	(fmap_rd_data_II[0]	),
    .\fmap_rd_data_II[1]	(fmap_rd_data_II[1]	),
    .\fmap_rd_data_II[2]	(fmap_rd_data_II[2]	),
    .\fmap_rd_data_II[3]	(fmap_rd_data_II[3]	),
    .\fmap_rd_data_II[4]	(fmap_rd_data_II[4]	),
    .\fmap_rd_data_II[5]	(fmap_rd_data_II[5]	),
    .\fmap_rd_data_II[6]	(fmap_rd_data_II[6]	),
    .\fmap_rd_data_II[7]	(fmap_rd_data_II[7]	),
    .\fmap_rd_data_II[8]	(fmap_rd_data_II[8]	),
    .\fmap_rd_data_II[9]	(fmap_rd_data_II[9]	),
    .\fmap_rd_data_II[10]	(fmap_rd_data_II[10]	),
    .\fmap_rd_data_II[11]	(fmap_rd_data_II[11]	),
    .\fmap_rd_data_II[12]	(fmap_rd_data_II[12]	),
    .\fmap_rd_data_II[13]	(fmap_rd_data_II[13]	),
    .\fmap_rd_data_II[14]	(fmap_rd_data_II[14]	),
    .\fmap_rd_data_II[15]	(fmap_rd_data_II[15]	),
    .\fmap_rd_data_II[16]	(fmap_rd_data_II[16]	),
    .\fmap_rd_data_II[17]	(fmap_rd_data_II[17]	),
    .\fmap_rd_data_II[18]	(fmap_rd_data_II[18]	),
    .\fmap_rd_data_II[19]	(fmap_rd_data_II[19]	),
    .\fmap_rd_data_II[20]	(fmap_rd_data_II[20]	),
    .\fmap_rd_data_II[21]	(fmap_rd_data_II[21]	),
    .\fmap_rd_data_II[22]	(fmap_rd_data_II[22]	),
    .\fmap_rd_data_II[23]	(fmap_rd_data_II[23]	),
    .\fmap_rd_data_II[24]	(fmap_rd_data_II[24]	),
    .\fmap_rd_data_II[25]	(fmap_rd_data_II[25]	),
    .\fmap_rd_data_II[26]	(fmap_rd_data_II[26]	),
    .\fmap_rd_data_II[27]	(fmap_rd_data_II[27]	),
    .\fmap_rd_data_II[28]	(fmap_rd_data_II[28]	),
    .\fmap_rd_data_II[29]	(fmap_rd_data_II[29]	),
    .\fmap_rd_data_II[30]	(fmap_rd_data_II[30]	),
    .\fmap_rd_data_II[31]	(fmap_rd_data_II[31]	),
    .\fmap_rd_data_II[32]	(fmap_rd_data_II[32]	),
    .\fmap_rd_data_II[33]	(fmap_rd_data_II[33]	),
    .\fmap_rd_data_II[34]	(fmap_rd_data_II[34]	),
    .\fmap_rd_data_II[35]	(fmap_rd_data_II[35]	),
    .\fmap_rd_data_II[36]	(fmap_rd_data_II[36]	),
    .\fmap_rd_data_II[37]	(fmap_rd_data_II[37]	),
    .\fmap_rd_data_II[38]	(fmap_rd_data_II[38]	),
    .\fmap_rd_data_II[39]	(fmap_rd_data_II[39]	),
    .\fmap_rd_data_II[40]	(fmap_rd_data_II[40]	),
    .\fmap_rd_data_II[41]	(fmap_rd_data_II[41]	),
    .\fmap_rd_data_II[42]	(fmap_rd_data_II[42]	),
    .\fmap_rd_data_II[43]	(fmap_rd_data_II[43]	),
    .\fmap_rd_data_II[44]	(fmap_rd_data_II[44]	),
    .\fmap_rd_data_II[45]	(fmap_rd_data_II[45]	),
    .\fmap_rd_data_II[46]	(fmap_rd_data_II[46]	),
    .\fmap_rd_data_II[47]	(fmap_rd_data_II[47]	),
    .\fmap_rd_data_II[48]	(fmap_rd_data_II[48]	),
    .\fmap_rd_data_II[49]	(fmap_rd_data_II[49]	),
    .\fmap_rd_data_II[50]	(fmap_rd_data_II[50]	),
    .\fmap_rd_data_II[51]	(fmap_rd_data_II[51]	),
    .\fmap_rd_data_II[52]	(fmap_rd_data_II[52]	),
    .\fmap_rd_data_II[53]	(fmap_rd_data_II[53]	),
    .\fmap_rd_data_II[54]	(fmap_rd_data_II[54]	),
    .\fmap_rd_data_II[55]	(fmap_rd_data_II[55]	),
    .\fmap_rd_data_II[56]	(fmap_rd_data_II[56]	),
    .\fmap_rd_data_II[57]	(fmap_rd_data_II[57]	),
    .\fmap_rd_data_II[58]	(fmap_rd_data_II[58]	),
    .\fmap_rd_data_II[59]	(fmap_rd_data_II[59]	),
    .\fmap_rd_data_II[60]	(fmap_rd_data_II[60]	),
    .\fmap_rd_data_II[61]	(fmap_rd_data_II[61]	),
    .\fmap_rd_data_II[62]	(fmap_rd_data_II[62]	),
    .\fmap_rd_data_II[63]	(fmap_rd_data_II[63]	),
    .\fmap_rd_data_II[64]	(fmap_rd_data_II[64]	),
    .\fmap_rd_data_II[65]	(fmap_rd_data_II[65]	),
    .\fmap_rd_data_II[66]	(fmap_rd_data_II[66]	),
    .\fmap_rd_data_II[67]	(fmap_rd_data_II[67]	),
    .\fmap_rd_data_II[68]	(fmap_rd_data_II[68]	),
    .\fmap_rd_data_II[69]	(fmap_rd_data_II[69]	),
    .\fmap_rd_data_II[70]	(fmap_rd_data_II[70]	),
    .\fmap_rd_data_II[71]	(fmap_rd_data_II[71]	),
    .\fmap_rd_data_II[72]	(fmap_rd_data_II[72]	),
    .\fmap_rd_data_II[73]	(fmap_rd_data_II[73]	),
    .\fmap_rd_data_II[74]	(fmap_rd_data_II[74]	),
    .\fmap_rd_data_II[75]	(fmap_rd_data_II[75]	),
    .\fmap_rd_data_II[76]	(fmap_rd_data_II[76]	),
    .\fmap_rd_data_II[77]	(fmap_rd_data_II[77]	),
    .\fmap_rd_data_II[78]	(fmap_rd_data_II[78]	),
    .\fmap_rd_data_II[79]	(fmap_rd_data_II[79]	),
    .\fmap_rd_data_II[80]	(fmap_rd_data_II[80]	),
    .\fmap_rd_data_II[81]	(fmap_rd_data_II[81]	),
    .\fmap_rd_data_II[82]	(fmap_rd_data_II[82]	),
    .\fmap_rd_data_II[83]	(fmap_rd_data_II[83]	),
    .\fmap_rd_data_II[84]	(fmap_rd_data_II[84]	),
    .\fmap_rd_data_II[85]	(fmap_rd_data_II[85]	),
    .\fmap_rd_data_II[86]	(fmap_rd_data_II[86]	),
    .\fmap_rd_data_II[87]	(fmap_rd_data_II[87]	),
    .\fmap_rd_data_II[88]	(fmap_rd_data_II[88]	),
    .\fmap_rd_data_II[89]	(fmap_rd_data_II[89]	),
    .\fmap_rd_data_II[90]	(fmap_rd_data_II[90]	),
    .\fmap_rd_data_II[91]	(fmap_rd_data_II[91]	),
    .\fmap_rd_data_II[92]	(fmap_rd_data_II[92]	),
    .\fmap_rd_data_II[93]	(fmap_rd_data_II[93]	),
    .\fmap_rd_data_II[94]	(fmap_rd_data_II[94]	),
    .\fmap_rd_data_II[95]	(fmap_rd_data_II[95]	),
    .\fmap_rd_data_II[96]	(fmap_rd_data_II[96]	),
    .\fmap_rd_data_II[97]	(fmap_rd_data_II[97]	),
    .\fmap_rd_data_II[98]	(fmap_rd_data_II[98]	),
    .\fmap_rd_data_II[99]	(fmap_rd_data_II[99]	),
    .\fmap_rd_data_II[100]	(fmap_rd_data_II[100]	),
    .\fmap_rd_data_II[101]	(fmap_rd_data_II[101]	),
    .\fmap_rd_data_II[102]	(fmap_rd_data_II[102]	),
    .\fmap_rd_data_II[103]	(fmap_rd_data_II[103]	),
    .\fmap_rd_data_II[104]	(fmap_rd_data_II[104]	),
    .\fmap_rd_data_II[105]	(fmap_rd_data_II[105]	),
    .\fmap_rd_data_II[106]	(fmap_rd_data_II[106]	),
    .\fmap_rd_data_II[107]	(fmap_rd_data_II[107]	),
    .\fmap_rd_data_II[108]	(fmap_rd_data_II[108]	),
    .\fmap_rd_data_II[109]	(fmap_rd_data_II[109]	),
    .\fmap_rd_data_II[110]	(fmap_rd_data_II[110]	),
    .\fmap_rd_data_II[111]	(fmap_rd_data_II[111]	),
    .\fmap_rd_data_II[112]	(fmap_rd_data_II[112]	),
    .\fmap_rd_data_II[113]	(fmap_rd_data_II[113]	),
    .\fmap_rd_data_II[114]	(fmap_rd_data_II[114]	),
    .\fmap_rd_data_II[115]	(fmap_rd_data_II[115]	),
    .\fmap_rd_data_II[116]	(fmap_rd_data_II[116]	),
    .\fmap_rd_data_II[117]	(fmap_rd_data_II[117]	),
    .\fmap_rd_data_II[118]	(fmap_rd_data_II[118]	),
    .\fmap_rd_data_II[119]	(fmap_rd_data_II[119]	),
    .\fmap_rd_data_II[120]	(fmap_rd_data_II[120]	),
    .\fmap_rd_data_II[121]	(fmap_rd_data_II[121]	),
    .\fmap_rd_data_II[122]	(fmap_rd_data_II[122]	),
    .\fmap_rd_data_II[123]	(fmap_rd_data_II[123]	),
    .\fmap_rd_data_II[124]	(fmap_rd_data_II[124]	),
    .\fmap_rd_data_II[125]	(fmap_rd_data_II[125]	),
    .\fmap_rd_data_II[126]	(fmap_rd_data_II[126]	),
    .\fmap_rd_data_II[127]	(fmap_rd_data_II[127]	),
    .\fmap_rd_data_II[128]	(fmap_rd_data_II[128]	),
    .\fmap_rd_data_II[129]	(fmap_rd_data_II[129]	),
    .\fmap_rd_data_II[130]	(fmap_rd_data_II[130]	),
    .\fmap_rd_data_II[131]	(fmap_rd_data_II[131]	),
    .\fmap_rd_data_II[132]	(fmap_rd_data_II[132]	),
    .\fmap_rd_data_II[133]	(fmap_rd_data_II[133]	),
    .\fmap_rd_data_II[134]	(fmap_rd_data_II[134]	),
    .\fmap_rd_data_II[135]	(fmap_rd_data_II[135]	),
    .\fmap_rd_data_II[136]	(fmap_rd_data_II[136]	),
    .\fmap_rd_data_II[137]	(fmap_rd_data_II[137]	),
    .\fmap_rd_data_II[138]	(fmap_rd_data_II[138]	),
    .\fmap_rd_data_II[139]	(fmap_rd_data_II[139]	),
    .\fmap_rd_data_II[140]	(fmap_rd_data_II[140]	),
    .\fmap_rd_data_II[141]	(fmap_rd_data_II[141]	),
    .\fmap_rd_data_II[142]	(fmap_rd_data_II[142]	),
    .\fmap_rd_data_II[143]	(fmap_rd_data_II[143]	),

    .\fmap_wr_data_II[0]	(fmap_wr_data_II[0]	),
    .\fmap_wr_data_II[1]	(fmap_wr_data_II[1]	),
    .\fmap_wr_data_II[2]	(fmap_wr_data_II[2]	),
    .\fmap_wr_data_II[3]	(fmap_wr_data_II[3]	),
    .\fmap_wr_data_II[4]	(fmap_wr_data_II[4]	),
    .\fmap_wr_data_II[5]	(fmap_wr_data_II[5]	),
    .\fmap_wr_data_II[6]	(fmap_wr_data_II[6]	),
    .\fmap_wr_data_II[7]	(fmap_wr_data_II[7]	),
    .\fmap_wr_data_II[8]	(fmap_wr_data_II[8]	),
    .\fmap_wr_data_II[9]	(fmap_wr_data_II[9]	),
    .\fmap_wr_data_II[10]	(fmap_wr_data_II[10]	),
    .\fmap_wr_data_II[11]	(fmap_wr_data_II[11]	),
    .\fmap_wr_data_II[12]	(fmap_wr_data_II[12]	),
    .\fmap_wr_data_II[13]	(fmap_wr_data_II[13]	),
    .\fmap_wr_data_II[14]	(fmap_wr_data_II[14]	),
    .\fmap_wr_data_II[15]	(fmap_wr_data_II[15]	),
    .\fmap_wr_data_II[16]	(fmap_wr_data_II[16]	),
    .\fmap_wr_data_II[17]	(fmap_wr_data_II[17]	),
    .\fmap_wr_data_II[18]	(fmap_wr_data_II[18]	),
    .\fmap_wr_data_II[19]	(fmap_wr_data_II[19]	),
    .\fmap_wr_data_II[20]	(fmap_wr_data_II[20]	),
    .\fmap_wr_data_II[21]	(fmap_wr_data_II[21]	),
    .\fmap_wr_data_II[22]	(fmap_wr_data_II[22]	),
    .\fmap_wr_data_II[23]	(fmap_wr_data_II[23]	),
    .\fmap_wr_data_II[24]	(fmap_wr_data_II[24]	),
    .\fmap_wr_data_II[25]	(fmap_wr_data_II[25]	),
    .\fmap_wr_data_II[26]	(fmap_wr_data_II[26]	),
    .\fmap_wr_data_II[27]	(fmap_wr_data_II[27]	),
    .\fmap_wr_data_II[28]	(fmap_wr_data_II[28]	),
    .\fmap_wr_data_II[29]	(fmap_wr_data_II[29]	),
    .\fmap_wr_data_II[30]	(fmap_wr_data_II[30]	),
    .\fmap_wr_data_II[31]	(fmap_wr_data_II[31]	),
    .\fmap_wr_data_II[32]	(fmap_wr_data_II[32]	),
    .\fmap_wr_data_II[33]	(fmap_wr_data_II[33]	),
    .\fmap_wr_data_II[34]	(fmap_wr_data_II[34]	),
    .\fmap_wr_data_II[35]	(fmap_wr_data_II[35]	),
    .\fmap_wr_data_II[36]	(fmap_wr_data_II[36]	),
    .\fmap_wr_data_II[37]	(fmap_wr_data_II[37]	),
    .\fmap_wr_data_II[38]	(fmap_wr_data_II[38]	),
    .\fmap_wr_data_II[39]	(fmap_wr_data_II[39]	),
    .\fmap_wr_data_II[40]	(fmap_wr_data_II[40]	),
    .\fmap_wr_data_II[41]	(fmap_wr_data_II[41]	),
    .\fmap_wr_data_II[42]	(fmap_wr_data_II[42]	),
    .\fmap_wr_data_II[43]	(fmap_wr_data_II[43]	),
    .\fmap_wr_data_II[44]	(fmap_wr_data_II[44]	),
    .\fmap_wr_data_II[45]	(fmap_wr_data_II[45]	),
    .\fmap_wr_data_II[46]	(fmap_wr_data_II[46]	),
    .\fmap_wr_data_II[47]	(fmap_wr_data_II[47]	),
    .\fmap_wr_data_II[48]	(fmap_wr_data_II[48]	),
    .\fmap_wr_data_II[49]	(fmap_wr_data_II[49]	),
    .\fmap_wr_data_II[50]	(fmap_wr_data_II[50]	),
    .\fmap_wr_data_II[51]	(fmap_wr_data_II[51]	),
    .\fmap_wr_data_II[52]	(fmap_wr_data_II[52]	),
    .\fmap_wr_data_II[53]	(fmap_wr_data_II[53]	),
    .\fmap_wr_data_II[54]	(fmap_wr_data_II[54]	),
    .\fmap_wr_data_II[55]	(fmap_wr_data_II[55]	),
    .\fmap_wr_data_II[56]	(fmap_wr_data_II[56]	),
    .\fmap_wr_data_II[57]	(fmap_wr_data_II[57]	),
    .\fmap_wr_data_II[58]	(fmap_wr_data_II[58]	),
    .\fmap_wr_data_II[59]	(fmap_wr_data_II[59]	),
    .\fmap_wr_data_II[60]	(fmap_wr_data_II[60]	),
    .\fmap_wr_data_II[61]	(fmap_wr_data_II[61]	),
    .\fmap_wr_data_II[62]	(fmap_wr_data_II[62]	),
    .\fmap_wr_data_II[63]	(fmap_wr_data_II[63]	),
    .\fmap_wr_data_II[64]	(fmap_wr_data_II[64]	),
    .\fmap_wr_data_II[65]	(fmap_wr_data_II[65]	),
    .\fmap_wr_data_II[66]	(fmap_wr_data_II[66]	),
    .\fmap_wr_data_II[67]	(fmap_wr_data_II[67]	),
    .\fmap_wr_data_II[68]	(fmap_wr_data_II[68]	),
    .\fmap_wr_data_II[69]	(fmap_wr_data_II[69]	),
    .\fmap_wr_data_II[70]	(fmap_wr_data_II[70]	),
    .\fmap_wr_data_II[71]	(fmap_wr_data_II[71]	),
    .\fmap_wr_data_II[72]	(fmap_wr_data_II[72]	),
    .\fmap_wr_data_II[73]	(fmap_wr_data_II[73]	),
    .\fmap_wr_data_II[74]	(fmap_wr_data_II[74]	),
    .\fmap_wr_data_II[75]	(fmap_wr_data_II[75]	),
    .\fmap_wr_data_II[76]	(fmap_wr_data_II[76]	),
    .\fmap_wr_data_II[77]	(fmap_wr_data_II[77]	),
    .\fmap_wr_data_II[78]	(fmap_wr_data_II[78]	),
    .\fmap_wr_data_II[79]	(fmap_wr_data_II[79]	),
    .\fmap_wr_data_II[80]	(fmap_wr_data_II[80]	),
    .\fmap_wr_data_II[81]	(fmap_wr_data_II[81]	),
    .\fmap_wr_data_II[82]	(fmap_wr_data_II[82]	),
    .\fmap_wr_data_II[83]	(fmap_wr_data_II[83]	),
    .\fmap_wr_data_II[84]	(fmap_wr_data_II[84]	),
    .\fmap_wr_data_II[85]	(fmap_wr_data_II[85]	),
    .\fmap_wr_data_II[86]	(fmap_wr_data_II[86]	),
    .\fmap_wr_data_II[87]	(fmap_wr_data_II[87]	),
    .\fmap_wr_data_II[88]	(fmap_wr_data_II[88]	),
    .\fmap_wr_data_II[89]	(fmap_wr_data_II[89]	),
    .\fmap_wr_data_II[90]	(fmap_wr_data_II[90]	),
    .\fmap_wr_data_II[91]	(fmap_wr_data_II[91]	),
    .\fmap_wr_data_II[92]	(fmap_wr_data_II[92]	),
    .\fmap_wr_data_II[93]	(fmap_wr_data_II[93]	),
    .\fmap_wr_data_II[94]	(fmap_wr_data_II[94]	),
    .\fmap_wr_data_II[95]	(fmap_wr_data_II[95]	),
    .\fmap_wr_data_II[96]	(fmap_wr_data_II[96]	),
    .\fmap_wr_data_II[97]	(fmap_wr_data_II[97]	),
    .\fmap_wr_data_II[98]	(fmap_wr_data_II[98]	),
    .\fmap_wr_data_II[99]	(fmap_wr_data_II[99]	),
    .\fmap_wr_data_II[100]	(fmap_wr_data_II[100]	),
    .\fmap_wr_data_II[101]	(fmap_wr_data_II[101]	),
    .\fmap_wr_data_II[102]	(fmap_wr_data_II[102]	),
    .\fmap_wr_data_II[103]	(fmap_wr_data_II[103]	),
    .\fmap_wr_data_II[104]	(fmap_wr_data_II[104]	),
    .\fmap_wr_data_II[105]	(fmap_wr_data_II[105]	),
    .\fmap_wr_data_II[106]	(fmap_wr_data_II[106]	),
    .\fmap_wr_data_II[107]	(fmap_wr_data_II[107]	),
    .\fmap_wr_data_II[108]	(fmap_wr_data_II[108]	),
    .\fmap_wr_data_II[109]	(fmap_wr_data_II[109]	),
    .\fmap_wr_data_II[110]	(fmap_wr_data_II[110]	),
    .\fmap_wr_data_II[111]	(fmap_wr_data_II[111]	),
    .\fmap_wr_data_II[112]	(fmap_wr_data_II[112]	),
    .\fmap_wr_data_II[113]	(fmap_wr_data_II[113]	),
    .\fmap_wr_data_II[114]	(fmap_wr_data_II[114]	),
    .\fmap_wr_data_II[115]	(fmap_wr_data_II[115]	),
    .\fmap_wr_data_II[116]	(fmap_wr_data_II[116]	),
    .\fmap_wr_data_II[117]	(fmap_wr_data_II[117]	),
    .\fmap_wr_data_II[118]	(fmap_wr_data_II[118]	),
    .\fmap_wr_data_II[119]	(fmap_wr_data_II[119]	),
    .\fmap_wr_data_II[120]	(fmap_wr_data_II[120]	),
    .\fmap_wr_data_II[121]	(fmap_wr_data_II[121]	),
    .\fmap_wr_data_II[122]	(fmap_wr_data_II[122]	),
    .\fmap_wr_data_II[123]	(fmap_wr_data_II[123]	),
    .\fmap_wr_data_II[124]	(fmap_wr_data_II[124]	),
    .\fmap_wr_data_II[125]	(fmap_wr_data_II[125]	),
    .\fmap_wr_data_II[126]	(fmap_wr_data_II[126]	),
    .\fmap_wr_data_II[127]	(fmap_wr_data_II[127]	),
    .\fmap_wr_data_II[128]	(fmap_wr_data_II[128]	),
    .\fmap_wr_data_II[129]	(fmap_wr_data_II[129]	),
    .\fmap_wr_data_II[130]	(fmap_wr_data_II[130]	),
    .\fmap_wr_data_II[131]	(fmap_wr_data_II[131]	),
    .\fmap_wr_data_II[132]	(fmap_wr_data_II[132]	),
    .\fmap_wr_data_II[133]	(fmap_wr_data_II[133]	),
    .\fmap_wr_data_II[134]	(fmap_wr_data_II[134]	),
    .\fmap_wr_data_II[135]	(fmap_wr_data_II[135]	),
    .\fmap_wr_data_II[136]	(fmap_wr_data_II[136]	),
    .\fmap_wr_data_II[137]	(fmap_wr_data_II[137]	),
    .\fmap_wr_data_II[138]	(fmap_wr_data_II[138]	),
    .\fmap_wr_data_II[139]	(fmap_wr_data_II[139]	),
    .\fmap_wr_data_II[140]	(fmap_wr_data_II[140]	),
    .\fmap_wr_data_II[141]	(fmap_wr_data_II[141]	),
    .\fmap_wr_data_II[142]	(fmap_wr_data_II[142]	),
    .\fmap_wr_data_II[143]	(fmap_wr_data_II[143]	),

    .\fmap_wr_en_II[0]	(fmap_wr_en_II[0]	),
    .\fmap_wr_en_II[1]	(fmap_wr_en_II[1]	),
    .\fmap_wr_en_II[2]	(fmap_wr_en_II[2]	),
    .\fmap_wr_en_II[3]	(fmap_wr_en_II[3]	),
    .\fmap_wr_en_II[4]	(fmap_wr_en_II[4]	),
    .\fmap_wr_en_II[5]	(fmap_wr_en_II[5]	),
    .\fmap_wr_en_II[6]	(fmap_wr_en_II[6]	),
    .\fmap_wr_en_II[7]	(fmap_wr_en_II[7]	),
    .\fmap_wr_en_II[8]	(fmap_wr_en_II[8]	),
    .\fmap_wr_en_II[9]	(fmap_wr_en_II[9]	),
    .\fmap_wr_en_II[10]	(fmap_wr_en_II[10]	),
    .\fmap_wr_en_II[11]	(fmap_wr_en_II[11]	),
    .\fmap_wr_en_II[12]	(fmap_wr_en_II[12]	),
    .\fmap_wr_en_II[13]	(fmap_wr_en_II[13]	),
    .\fmap_wr_en_II[14]	(fmap_wr_en_II[14]	),
    .\fmap_wr_en_II[15]	(fmap_wr_en_II[15]	),
    .\fmap_wr_en_II[16]	(fmap_wr_en_II[16]	),
    .\fmap_wr_en_II[17]	(fmap_wr_en_II[17]	),
    .\fmap_wr_en_II[18]	(fmap_wr_en_II[18]	),
    .\fmap_wr_en_II[19]	(fmap_wr_en_II[19]	),
    .\fmap_wr_en_II[20]	(fmap_wr_en_II[20]	),
    .\fmap_wr_en_II[21]	(fmap_wr_en_II[21]	),
    .\fmap_wr_en_II[22]	(fmap_wr_en_II[22]	),
    .\fmap_wr_en_II[23]	(fmap_wr_en_II[23]	),
    .\fmap_wr_en_II[24]	(fmap_wr_en_II[24]	),
    .\fmap_wr_en_II[25]	(fmap_wr_en_II[25]	),
    .\fmap_wr_en_II[26]	(fmap_wr_en_II[26]	),
    .\fmap_wr_en_II[27]	(fmap_wr_en_II[27]	),
    .\fmap_wr_en_II[28]	(fmap_wr_en_II[28]	),
    .\fmap_wr_en_II[29]	(fmap_wr_en_II[29]	),
    .\fmap_wr_en_II[30]	(fmap_wr_en_II[30]	),
    .\fmap_wr_en_II[31]	(fmap_wr_en_II[31]	),
    .\fmap_wr_en_II[32]	(fmap_wr_en_II[32]	),
    .\fmap_wr_en_II[33]	(fmap_wr_en_II[33]	),
    .\fmap_wr_en_II[34]	(fmap_wr_en_II[34]	),
    .\fmap_wr_en_II[35]	(fmap_wr_en_II[35]	),
    .\fmap_wr_en_II[36]	(fmap_wr_en_II[36]	),
    .\fmap_wr_en_II[37]	(fmap_wr_en_II[37]	),
    .\fmap_wr_en_II[38]	(fmap_wr_en_II[38]	),
    .\fmap_wr_en_II[39]	(fmap_wr_en_II[39]	),
    .\fmap_wr_en_II[40]	(fmap_wr_en_II[40]	),
    .\fmap_wr_en_II[41]	(fmap_wr_en_II[41]	),
    .\fmap_wr_en_II[42]	(fmap_wr_en_II[42]	),
    .\fmap_wr_en_II[43]	(fmap_wr_en_II[43]	),
    .\fmap_wr_en_II[44]	(fmap_wr_en_II[44]	),
    .\fmap_wr_en_II[45]	(fmap_wr_en_II[45]	),
    .\fmap_wr_en_II[46]	(fmap_wr_en_II[46]	),
    .\fmap_wr_en_II[47]	(fmap_wr_en_II[47]	),
    .\fmap_wr_en_II[48]	(fmap_wr_en_II[48]	),
    .\fmap_wr_en_II[49]	(fmap_wr_en_II[49]	),
    .\fmap_wr_en_II[50]	(fmap_wr_en_II[50]	),
    .\fmap_wr_en_II[51]	(fmap_wr_en_II[51]	),
    .\fmap_wr_en_II[52]	(fmap_wr_en_II[52]	),
    .\fmap_wr_en_II[53]	(fmap_wr_en_II[53]	),
    .\fmap_wr_en_II[54]	(fmap_wr_en_II[54]	),
    .\fmap_wr_en_II[55]	(fmap_wr_en_II[55]	),
    .\fmap_wr_en_II[56]	(fmap_wr_en_II[56]	),
    .\fmap_wr_en_II[57]	(fmap_wr_en_II[57]	),
    .\fmap_wr_en_II[58]	(fmap_wr_en_II[58]	),
    .\fmap_wr_en_II[59]	(fmap_wr_en_II[59]	),
    .\fmap_wr_en_II[60]	(fmap_wr_en_II[60]	),
    .\fmap_wr_en_II[61]	(fmap_wr_en_II[61]	),
    .\fmap_wr_en_II[62]	(fmap_wr_en_II[62]	),
    .\fmap_wr_en_II[63]	(fmap_wr_en_II[63]	),
    .\fmap_wr_en_II[64]	(fmap_wr_en_II[64]	),
    .\fmap_wr_en_II[65]	(fmap_wr_en_II[65]	),
    .\fmap_wr_en_II[66]	(fmap_wr_en_II[66]	),
    .\fmap_wr_en_II[67]	(fmap_wr_en_II[67]	),
    .\fmap_wr_en_II[68]	(fmap_wr_en_II[68]	),
    .\fmap_wr_en_II[69]	(fmap_wr_en_II[69]	),
    .\fmap_wr_en_II[70]	(fmap_wr_en_II[70]	),
    .\fmap_wr_en_II[71]	(fmap_wr_en_II[71]	),
    .\fmap_wr_en_II[72]	(fmap_wr_en_II[72]	),
    .\fmap_wr_en_II[73]	(fmap_wr_en_II[73]	),
    .\fmap_wr_en_II[74]	(fmap_wr_en_II[74]	),
    .\fmap_wr_en_II[75]	(fmap_wr_en_II[75]	),
    .\fmap_wr_en_II[76]	(fmap_wr_en_II[76]	),
    .\fmap_wr_en_II[77]	(fmap_wr_en_II[77]	),
    .\fmap_wr_en_II[78]	(fmap_wr_en_II[78]	),
    .\fmap_wr_en_II[79]	(fmap_wr_en_II[79]	),
    .\fmap_wr_en_II[80]	(fmap_wr_en_II[80]	),
    .\fmap_wr_en_II[81]	(fmap_wr_en_II[81]	),
    .\fmap_wr_en_II[82]	(fmap_wr_en_II[82]	),
    .\fmap_wr_en_II[83]	(fmap_wr_en_II[83]	),
    .\fmap_wr_en_II[84]	(fmap_wr_en_II[84]	),
    .\fmap_wr_en_II[85]	(fmap_wr_en_II[85]	),
    .\fmap_wr_en_II[86]	(fmap_wr_en_II[86]	),
    .\fmap_wr_en_II[87]	(fmap_wr_en_II[87]	),
    .\fmap_wr_en_II[88]	(fmap_wr_en_II[88]	),
    .\fmap_wr_en_II[89]	(fmap_wr_en_II[89]	),
    .\fmap_wr_en_II[90]	(fmap_wr_en_II[90]	),
    .\fmap_wr_en_II[91]	(fmap_wr_en_II[91]	),
    .\fmap_wr_en_II[92]	(fmap_wr_en_II[92]	),
    .\fmap_wr_en_II[93]	(fmap_wr_en_II[93]	),
    .\fmap_wr_en_II[94]	(fmap_wr_en_II[94]	),
    .\fmap_wr_en_II[95]	(fmap_wr_en_II[95]	),
    .\fmap_wr_en_II[96]	(fmap_wr_en_II[96]	),
    .\fmap_wr_en_II[97]	(fmap_wr_en_II[97]	),
    .\fmap_wr_en_II[98]	(fmap_wr_en_II[98]	),
    .\fmap_wr_en_II[99]	(fmap_wr_en_II[99]	),
    .\fmap_wr_en_II[100]	(fmap_wr_en_II[100]	),
    .\fmap_wr_en_II[101]	(fmap_wr_en_II[101]	),
    .\fmap_wr_en_II[102]	(fmap_wr_en_II[102]	),
    .\fmap_wr_en_II[103]	(fmap_wr_en_II[103]	),
    .\fmap_wr_en_II[104]	(fmap_wr_en_II[104]	),
    .\fmap_wr_en_II[105]	(fmap_wr_en_II[105]	),
    .\fmap_wr_en_II[106]	(fmap_wr_en_II[106]	),
    .\fmap_wr_en_II[107]	(fmap_wr_en_II[107]	),
    .\fmap_wr_en_II[108]	(fmap_wr_en_II[108]	),
    .\fmap_wr_en_II[109]	(fmap_wr_en_II[109]	),
    .\fmap_wr_en_II[110]	(fmap_wr_en_II[110]	),
    .\fmap_wr_en_II[111]	(fmap_wr_en_II[111]	),
    .\fmap_wr_en_II[112]	(fmap_wr_en_II[112]	),
    .\fmap_wr_en_II[113]	(fmap_wr_en_II[113]	),
    .\fmap_wr_en_II[114]	(fmap_wr_en_II[114]	),
    .\fmap_wr_en_II[115]	(fmap_wr_en_II[115]	),
    .\fmap_wr_en_II[116]	(fmap_wr_en_II[116]	),
    .\fmap_wr_en_II[117]	(fmap_wr_en_II[117]	),
    .\fmap_wr_en_II[118]	(fmap_wr_en_II[118]	),
    .\fmap_wr_en_II[119]	(fmap_wr_en_II[119]	),
    .\fmap_wr_en_II[120]	(fmap_wr_en_II[120]	),
    .\fmap_wr_en_II[121]	(fmap_wr_en_II[121]	),
    .\fmap_wr_en_II[122]	(fmap_wr_en_II[122]	),
    .\fmap_wr_en_II[123]	(fmap_wr_en_II[123]	),
    .\fmap_wr_en_II[124]	(fmap_wr_en_II[124]	),
    .\fmap_wr_en_II[125]	(fmap_wr_en_II[125]	),
    .\fmap_wr_en_II[126]	(fmap_wr_en_II[126]	),
    .\fmap_wr_en_II[127]	(fmap_wr_en_II[127]	),
    .\fmap_wr_en_II[128]	(fmap_wr_en_II[128]	),
    .\fmap_wr_en_II[129]	(fmap_wr_en_II[129]	),
    .\fmap_wr_en_II[130]	(fmap_wr_en_II[130]	),
    .\fmap_wr_en_II[131]	(fmap_wr_en_II[131]	),
    .\fmap_wr_en_II[132]	(fmap_wr_en_II[132]	),
    .\fmap_wr_en_II[133]	(fmap_wr_en_II[133]	),
    .\fmap_wr_en_II[134]	(fmap_wr_en_II[134]	),
    .\fmap_wr_en_II[135]	(fmap_wr_en_II[135]	),
    .\fmap_wr_en_II[136]	(fmap_wr_en_II[136]	),
    .\fmap_wr_en_II[137]	(fmap_wr_en_II[137]	),
    .\fmap_wr_en_II[138]	(fmap_wr_en_II[138]	),
    .\fmap_wr_en_II[139]	(fmap_wr_en_II[139]	),
    .\fmap_wr_en_II[140]	(fmap_wr_en_II[140]	),
    .\fmap_wr_en_II[141]	(fmap_wr_en_II[141]	),
    .\fmap_wr_en_II[142]	(fmap_wr_en_II[142]	),
    .\fmap_wr_en_II[143]	(fmap_wr_en_II[143]	),

    .\fmap_wr_addr_II[0]	(fmap_wr_addr_II[0]	),
    .\fmap_wr_addr_II[1]	(fmap_wr_addr_II[1]	),
    .\fmap_wr_addr_II[2]	(fmap_wr_addr_II[2]	),
    .\fmap_wr_addr_II[3]	(fmap_wr_addr_II[3]	),
    .\fmap_wr_addr_II[4]	(fmap_wr_addr_II[4]	),
    .\fmap_wr_addr_II[5]	(fmap_wr_addr_II[5]	),
    .\fmap_wr_addr_II[6]	(fmap_wr_addr_II[6]	),
    .\fmap_wr_addr_II[7]	(fmap_wr_addr_II[7]	),
    .\fmap_wr_addr_II[8]	(fmap_wr_addr_II[8]	),
    .\fmap_wr_addr_II[9]	(fmap_wr_addr_II[9]	),
    .\fmap_wr_addr_II[10]	(fmap_wr_addr_II[10]	),
    .\fmap_wr_addr_II[11]	(fmap_wr_addr_II[11]	),
    .\fmap_wr_addr_II[12]	(fmap_wr_addr_II[12]	),
    .\fmap_wr_addr_II[13]	(fmap_wr_addr_II[13]	),
    .\fmap_wr_addr_II[14]	(fmap_wr_addr_II[14]	),
    .\fmap_wr_addr_II[15]	(fmap_wr_addr_II[15]	),
    .\fmap_wr_addr_II[16]	(fmap_wr_addr_II[16]	),
    .\fmap_wr_addr_II[17]	(fmap_wr_addr_II[17]	),
    .\fmap_wr_addr_II[18]	(fmap_wr_addr_II[18]	),
    .\fmap_wr_addr_II[19]	(fmap_wr_addr_II[19]	),
    .\fmap_wr_addr_II[20]	(fmap_wr_addr_II[20]	),
    .\fmap_wr_addr_II[21]	(fmap_wr_addr_II[21]	),
    .\fmap_wr_addr_II[22]	(fmap_wr_addr_II[22]	),
    .\fmap_wr_addr_II[23]	(fmap_wr_addr_II[23]	),
    .\fmap_wr_addr_II[24]	(fmap_wr_addr_II[24]	),
    .\fmap_wr_addr_II[25]	(fmap_wr_addr_II[25]	),
    .\fmap_wr_addr_II[26]	(fmap_wr_addr_II[26]	),
    .\fmap_wr_addr_II[27]	(fmap_wr_addr_II[27]	),
    .\fmap_wr_addr_II[28]	(fmap_wr_addr_II[28]	),
    .\fmap_wr_addr_II[29]	(fmap_wr_addr_II[29]	),
    .\fmap_wr_addr_II[30]	(fmap_wr_addr_II[30]	),
    .\fmap_wr_addr_II[31]	(fmap_wr_addr_II[31]	),
    .\fmap_wr_addr_II[32]	(fmap_wr_addr_II[32]	),
    .\fmap_wr_addr_II[33]	(fmap_wr_addr_II[33]	),
    .\fmap_wr_addr_II[34]	(fmap_wr_addr_II[34]	),
    .\fmap_wr_addr_II[35]	(fmap_wr_addr_II[35]	),
    .\fmap_wr_addr_II[36]	(fmap_wr_addr_II[36]	),
    .\fmap_wr_addr_II[37]	(fmap_wr_addr_II[37]	),
    .\fmap_wr_addr_II[38]	(fmap_wr_addr_II[38]	),
    .\fmap_wr_addr_II[39]	(fmap_wr_addr_II[39]	),
    .\fmap_wr_addr_II[40]	(fmap_wr_addr_II[40]	),
    .\fmap_wr_addr_II[41]	(fmap_wr_addr_II[41]	),
    .\fmap_wr_addr_II[42]	(fmap_wr_addr_II[42]	),
    .\fmap_wr_addr_II[43]	(fmap_wr_addr_II[43]	),
    .\fmap_wr_addr_II[44]	(fmap_wr_addr_II[44]	),
    .\fmap_wr_addr_II[45]	(fmap_wr_addr_II[45]	),
    .\fmap_wr_addr_II[46]	(fmap_wr_addr_II[46]	),
    .\fmap_wr_addr_II[47]	(fmap_wr_addr_II[47]	),
    .\fmap_wr_addr_II[48]	(fmap_wr_addr_II[48]	),
    .\fmap_wr_addr_II[49]	(fmap_wr_addr_II[49]	),
    .\fmap_wr_addr_II[50]	(fmap_wr_addr_II[50]	),
    .\fmap_wr_addr_II[51]	(fmap_wr_addr_II[51]	),
    .\fmap_wr_addr_II[52]	(fmap_wr_addr_II[52]	),
    .\fmap_wr_addr_II[53]	(fmap_wr_addr_II[53]	),
    .\fmap_wr_addr_II[54]	(fmap_wr_addr_II[54]	),
    .\fmap_wr_addr_II[55]	(fmap_wr_addr_II[55]	),
    .\fmap_wr_addr_II[56]	(fmap_wr_addr_II[56]	),
    .\fmap_wr_addr_II[57]	(fmap_wr_addr_II[57]	),
    .\fmap_wr_addr_II[58]	(fmap_wr_addr_II[58]	),
    .\fmap_wr_addr_II[59]	(fmap_wr_addr_II[59]	),
    .\fmap_wr_addr_II[60]	(fmap_wr_addr_II[60]	),
    .\fmap_wr_addr_II[61]	(fmap_wr_addr_II[61]	),
    .\fmap_wr_addr_II[62]	(fmap_wr_addr_II[62]	),
    .\fmap_wr_addr_II[63]	(fmap_wr_addr_II[63]	),
    .\fmap_wr_addr_II[64]	(fmap_wr_addr_II[64]	),
    .\fmap_wr_addr_II[65]	(fmap_wr_addr_II[65]	),
    .\fmap_wr_addr_II[66]	(fmap_wr_addr_II[66]	),
    .\fmap_wr_addr_II[67]	(fmap_wr_addr_II[67]	),
    .\fmap_wr_addr_II[68]	(fmap_wr_addr_II[68]	),
    .\fmap_wr_addr_II[69]	(fmap_wr_addr_II[69]	),
    .\fmap_wr_addr_II[70]	(fmap_wr_addr_II[70]	),
    .\fmap_wr_addr_II[71]	(fmap_wr_addr_II[71]	),
    .\fmap_wr_addr_II[72]	(fmap_wr_addr_II[72]	),
    .\fmap_wr_addr_II[73]	(fmap_wr_addr_II[73]	),
    .\fmap_wr_addr_II[74]	(fmap_wr_addr_II[74]	),
    .\fmap_wr_addr_II[75]	(fmap_wr_addr_II[75]	),
    .\fmap_wr_addr_II[76]	(fmap_wr_addr_II[76]	),
    .\fmap_wr_addr_II[77]	(fmap_wr_addr_II[77]	),
    .\fmap_wr_addr_II[78]	(fmap_wr_addr_II[78]	),
    .\fmap_wr_addr_II[79]	(fmap_wr_addr_II[79]	),
    .\fmap_wr_addr_II[80]	(fmap_wr_addr_II[80]	),
    .\fmap_wr_addr_II[81]	(fmap_wr_addr_II[81]	),
    .\fmap_wr_addr_II[82]	(fmap_wr_addr_II[82]	),
    .\fmap_wr_addr_II[83]	(fmap_wr_addr_II[83]	),
    .\fmap_wr_addr_II[84]	(fmap_wr_addr_II[84]	),
    .\fmap_wr_addr_II[85]	(fmap_wr_addr_II[85]	),
    .\fmap_wr_addr_II[86]	(fmap_wr_addr_II[86]	),
    .\fmap_wr_addr_II[87]	(fmap_wr_addr_II[87]	),
    .\fmap_wr_addr_II[88]	(fmap_wr_addr_II[88]	),
    .\fmap_wr_addr_II[89]	(fmap_wr_addr_II[89]	),
    .\fmap_wr_addr_II[90]	(fmap_wr_addr_II[90]	),
    .\fmap_wr_addr_II[91]	(fmap_wr_addr_II[91]	),
    .\fmap_wr_addr_II[92]	(fmap_wr_addr_II[92]	),
    .\fmap_wr_addr_II[93]	(fmap_wr_addr_II[93]	),
    .\fmap_wr_addr_II[94]	(fmap_wr_addr_II[94]	),
    .\fmap_wr_addr_II[95]	(fmap_wr_addr_II[95]	),
    .\fmap_wr_addr_II[96]	(fmap_wr_addr_II[96]	),
    .\fmap_wr_addr_II[97]	(fmap_wr_addr_II[97]	),
    .\fmap_wr_addr_II[98]	(fmap_wr_addr_II[98]	),
    .\fmap_wr_addr_II[99]	(fmap_wr_addr_II[99]	),
    .\fmap_wr_addr_II[100]	(fmap_wr_addr_II[100]	),
    .\fmap_wr_addr_II[101]	(fmap_wr_addr_II[101]	),
    .\fmap_wr_addr_II[102]	(fmap_wr_addr_II[102]	),
    .\fmap_wr_addr_II[103]	(fmap_wr_addr_II[103]	),
    .\fmap_wr_addr_II[104]	(fmap_wr_addr_II[104]	),
    .\fmap_wr_addr_II[105]	(fmap_wr_addr_II[105]	),
    .\fmap_wr_addr_II[106]	(fmap_wr_addr_II[106]	),
    .\fmap_wr_addr_II[107]	(fmap_wr_addr_II[107]	),
    .\fmap_wr_addr_II[108]	(fmap_wr_addr_II[108]	),
    .\fmap_wr_addr_II[109]	(fmap_wr_addr_II[109]	),
    .\fmap_wr_addr_II[110]	(fmap_wr_addr_II[110]	),
    .\fmap_wr_addr_II[111]	(fmap_wr_addr_II[111]	),
    .\fmap_wr_addr_II[112]	(fmap_wr_addr_II[112]	),
    .\fmap_wr_addr_II[113]	(fmap_wr_addr_II[113]	),
    .\fmap_wr_addr_II[114]	(fmap_wr_addr_II[114]	),
    .\fmap_wr_addr_II[115]	(fmap_wr_addr_II[115]	),
    .\fmap_wr_addr_II[116]	(fmap_wr_addr_II[116]	),
    .\fmap_wr_addr_II[117]	(fmap_wr_addr_II[117]	),
    .\fmap_wr_addr_II[118]	(fmap_wr_addr_II[118]	),
    .\fmap_wr_addr_II[119]	(fmap_wr_addr_II[119]	),
    .\fmap_wr_addr_II[120]	(fmap_wr_addr_II[120]	),
    .\fmap_wr_addr_II[121]	(fmap_wr_addr_II[121]	),
    .\fmap_wr_addr_II[122]	(fmap_wr_addr_II[122]	),
    .\fmap_wr_addr_II[123]	(fmap_wr_addr_II[123]	),
    .\fmap_wr_addr_II[124]	(fmap_wr_addr_II[124]	),
    .\fmap_wr_addr_II[125]	(fmap_wr_addr_II[125]	),
    .\fmap_wr_addr_II[126]	(fmap_wr_addr_II[126]	),
    .\fmap_wr_addr_II[127]	(fmap_wr_addr_II[127]	),
    .\fmap_wr_addr_II[128]	(fmap_wr_addr_II[128]	),
    .\fmap_wr_addr_II[129]	(fmap_wr_addr_II[129]	),
    .\fmap_wr_addr_II[130]	(fmap_wr_addr_II[130]	),
    .\fmap_wr_addr_II[131]	(fmap_wr_addr_II[131]	),
    .\fmap_wr_addr_II[132]	(fmap_wr_addr_II[132]	),
    .\fmap_wr_addr_II[133]	(fmap_wr_addr_II[133]	),
    .\fmap_wr_addr_II[134]	(fmap_wr_addr_II[134]	),
    .\fmap_wr_addr_II[135]	(fmap_wr_addr_II[135]	),
    .\fmap_wr_addr_II[136]	(fmap_wr_addr_II[136]	),
    .\fmap_wr_addr_II[137]	(fmap_wr_addr_II[137]	),
    .\fmap_wr_addr_II[138]	(fmap_wr_addr_II[138]	),
    .\fmap_wr_addr_II[139]	(fmap_wr_addr_II[139]	),
    .\fmap_wr_addr_II[140]	(fmap_wr_addr_II[140]	),
    .\fmap_wr_addr_II[141]	(fmap_wr_addr_II[141]	),
    .\fmap_wr_addr_II[142]	(fmap_wr_addr_II[142]	),
    .\fmap_wr_addr_II[143]	(fmap_wr_addr_II[143]	),

    .\fmap_rd_addr_II[0]	(fmap_rd_addr_II[0]	),
    .\fmap_rd_addr_II[1]	(fmap_rd_addr_II[1]	),
    .\fmap_rd_addr_II[2]	(fmap_rd_addr_II[2]	),
    .\fmap_rd_addr_II[3]	(fmap_rd_addr_II[3]	),
    .\fmap_rd_addr_II[4]	(fmap_rd_addr_II[4]	),
    .\fmap_rd_addr_II[5]	(fmap_rd_addr_II[5]	),
    .\fmap_rd_addr_II[6]	(fmap_rd_addr_II[6]	),
    .\fmap_rd_addr_II[7]	(fmap_rd_addr_II[7]	),
    .\fmap_rd_addr_II[8]	(fmap_rd_addr_II[8]	),
    .\fmap_rd_addr_II[9]	(fmap_rd_addr_II[9]	),
    .\fmap_rd_addr_II[10]	(fmap_rd_addr_II[10]	),
    .\fmap_rd_addr_II[11]	(fmap_rd_addr_II[11]	),
    .\fmap_rd_addr_II[12]	(fmap_rd_addr_II[12]	),
    .\fmap_rd_addr_II[13]	(fmap_rd_addr_II[13]	),
    .\fmap_rd_addr_II[14]	(fmap_rd_addr_II[14]	),
    .\fmap_rd_addr_II[15]	(fmap_rd_addr_II[15]	),
    .\fmap_rd_addr_II[16]	(fmap_rd_addr_II[16]	),
    .\fmap_rd_addr_II[17]	(fmap_rd_addr_II[17]	),
    .\fmap_rd_addr_II[18]	(fmap_rd_addr_II[18]	),
    .\fmap_rd_addr_II[19]	(fmap_rd_addr_II[19]	),
    .\fmap_rd_addr_II[20]	(fmap_rd_addr_II[20]	),
    .\fmap_rd_addr_II[21]	(fmap_rd_addr_II[21]	),
    .\fmap_rd_addr_II[22]	(fmap_rd_addr_II[22]	),
    .\fmap_rd_addr_II[23]	(fmap_rd_addr_II[23]	),
    .\fmap_rd_addr_II[24]	(fmap_rd_addr_II[24]	),
    .\fmap_rd_addr_II[25]	(fmap_rd_addr_II[25]	),
    .\fmap_rd_addr_II[26]	(fmap_rd_addr_II[26]	),
    .\fmap_rd_addr_II[27]	(fmap_rd_addr_II[27]	),
    .\fmap_rd_addr_II[28]	(fmap_rd_addr_II[28]	),
    .\fmap_rd_addr_II[29]	(fmap_rd_addr_II[29]	),
    .\fmap_rd_addr_II[30]	(fmap_rd_addr_II[30]	),
    .\fmap_rd_addr_II[31]	(fmap_rd_addr_II[31]	),
    .\fmap_rd_addr_II[32]	(fmap_rd_addr_II[32]	),
    .\fmap_rd_addr_II[33]	(fmap_rd_addr_II[33]	),
    .\fmap_rd_addr_II[34]	(fmap_rd_addr_II[34]	),
    .\fmap_rd_addr_II[35]	(fmap_rd_addr_II[35]	),
    .\fmap_rd_addr_II[36]	(fmap_rd_addr_II[36]	),
    .\fmap_rd_addr_II[37]	(fmap_rd_addr_II[37]	),
    .\fmap_rd_addr_II[38]	(fmap_rd_addr_II[38]	),
    .\fmap_rd_addr_II[39]	(fmap_rd_addr_II[39]	),
    .\fmap_rd_addr_II[40]	(fmap_rd_addr_II[40]	),
    .\fmap_rd_addr_II[41]	(fmap_rd_addr_II[41]	),
    .\fmap_rd_addr_II[42]	(fmap_rd_addr_II[42]	),
    .\fmap_rd_addr_II[43]	(fmap_rd_addr_II[43]	),
    .\fmap_rd_addr_II[44]	(fmap_rd_addr_II[44]	),
    .\fmap_rd_addr_II[45]	(fmap_rd_addr_II[45]	),
    .\fmap_rd_addr_II[46]	(fmap_rd_addr_II[46]	),
    .\fmap_rd_addr_II[47]	(fmap_rd_addr_II[47]	),
    .\fmap_rd_addr_II[48]	(fmap_rd_addr_II[48]	),
    .\fmap_rd_addr_II[49]	(fmap_rd_addr_II[49]	),
    .\fmap_rd_addr_II[50]	(fmap_rd_addr_II[50]	),
    .\fmap_rd_addr_II[51]	(fmap_rd_addr_II[51]	),
    .\fmap_rd_addr_II[52]	(fmap_rd_addr_II[52]	),
    .\fmap_rd_addr_II[53]	(fmap_rd_addr_II[53]	),
    .\fmap_rd_addr_II[54]	(fmap_rd_addr_II[54]	),
    .\fmap_rd_addr_II[55]	(fmap_rd_addr_II[55]	),
    .\fmap_rd_addr_II[56]	(fmap_rd_addr_II[56]	),
    .\fmap_rd_addr_II[57]	(fmap_rd_addr_II[57]	),
    .\fmap_rd_addr_II[58]	(fmap_rd_addr_II[58]	),
    .\fmap_rd_addr_II[59]	(fmap_rd_addr_II[59]	),
    .\fmap_rd_addr_II[60]	(fmap_rd_addr_II[60]	),
    .\fmap_rd_addr_II[61]	(fmap_rd_addr_II[61]	),
    .\fmap_rd_addr_II[62]	(fmap_rd_addr_II[62]	),
    .\fmap_rd_addr_II[63]	(fmap_rd_addr_II[63]	),
    .\fmap_rd_addr_II[64]	(fmap_rd_addr_II[64]	),
    .\fmap_rd_addr_II[65]	(fmap_rd_addr_II[65]	),
    .\fmap_rd_addr_II[66]	(fmap_rd_addr_II[66]	),
    .\fmap_rd_addr_II[67]	(fmap_rd_addr_II[67]	),
    .\fmap_rd_addr_II[68]	(fmap_rd_addr_II[68]	),
    .\fmap_rd_addr_II[69]	(fmap_rd_addr_II[69]	),
    .\fmap_rd_addr_II[70]	(fmap_rd_addr_II[70]	),
    .\fmap_rd_addr_II[71]	(fmap_rd_addr_II[71]	),
    .\fmap_rd_addr_II[72]	(fmap_rd_addr_II[72]	),
    .\fmap_rd_addr_II[73]	(fmap_rd_addr_II[73]	),
    .\fmap_rd_addr_II[74]	(fmap_rd_addr_II[74]	),
    .\fmap_rd_addr_II[75]	(fmap_rd_addr_II[75]	),
    .\fmap_rd_addr_II[76]	(fmap_rd_addr_II[76]	),
    .\fmap_rd_addr_II[77]	(fmap_rd_addr_II[77]	),
    .\fmap_rd_addr_II[78]	(fmap_rd_addr_II[78]	),
    .\fmap_rd_addr_II[79]	(fmap_rd_addr_II[79]	),
    .\fmap_rd_addr_II[80]	(fmap_rd_addr_II[80]	),
    .\fmap_rd_addr_II[81]	(fmap_rd_addr_II[81]	),
    .\fmap_rd_addr_II[82]	(fmap_rd_addr_II[82]	),
    .\fmap_rd_addr_II[83]	(fmap_rd_addr_II[83]	),
    .\fmap_rd_addr_II[84]	(fmap_rd_addr_II[84]	),
    .\fmap_rd_addr_II[85]	(fmap_rd_addr_II[85]	),
    .\fmap_rd_addr_II[86]	(fmap_rd_addr_II[86]	),
    .\fmap_rd_addr_II[87]	(fmap_rd_addr_II[87]	),
    .\fmap_rd_addr_II[88]	(fmap_rd_addr_II[88]	),
    .\fmap_rd_addr_II[89]	(fmap_rd_addr_II[89]	),
    .\fmap_rd_addr_II[90]	(fmap_rd_addr_II[90]	),
    .\fmap_rd_addr_II[91]	(fmap_rd_addr_II[91]	),
    .\fmap_rd_addr_II[92]	(fmap_rd_addr_II[92]	),
    .\fmap_rd_addr_II[93]	(fmap_rd_addr_II[93]	),
    .\fmap_rd_addr_II[94]	(fmap_rd_addr_II[94]	),
    .\fmap_rd_addr_II[95]	(fmap_rd_addr_II[95]	),
    .\fmap_rd_addr_II[96]	(fmap_rd_addr_II[96]	),
    .\fmap_rd_addr_II[97]	(fmap_rd_addr_II[97]	),
    .\fmap_rd_addr_II[98]	(fmap_rd_addr_II[98]	),
    .\fmap_rd_addr_II[99]	(fmap_rd_addr_II[99]	),
    .\fmap_rd_addr_II[100]	(fmap_rd_addr_II[100]	),
    .\fmap_rd_addr_II[101]	(fmap_rd_addr_II[101]	),
    .\fmap_rd_addr_II[102]	(fmap_rd_addr_II[102]	),
    .\fmap_rd_addr_II[103]	(fmap_rd_addr_II[103]	),
    .\fmap_rd_addr_II[104]	(fmap_rd_addr_II[104]	),
    .\fmap_rd_addr_II[105]	(fmap_rd_addr_II[105]	),
    .\fmap_rd_addr_II[106]	(fmap_rd_addr_II[106]	),
    .\fmap_rd_addr_II[107]	(fmap_rd_addr_II[107]	),
    .\fmap_rd_addr_II[108]	(fmap_rd_addr_II[108]	),
    .\fmap_rd_addr_II[109]	(fmap_rd_addr_II[109]	),
    .\fmap_rd_addr_II[110]	(fmap_rd_addr_II[110]	),
    .\fmap_rd_addr_II[111]	(fmap_rd_addr_II[111]	),
    .\fmap_rd_addr_II[112]	(fmap_rd_addr_II[112]	),
    .\fmap_rd_addr_II[113]	(fmap_rd_addr_II[113]	),
    .\fmap_rd_addr_II[114]	(fmap_rd_addr_II[114]	),
    .\fmap_rd_addr_II[115]	(fmap_rd_addr_II[115]	),
    .\fmap_rd_addr_II[116]	(fmap_rd_addr_II[116]	),
    .\fmap_rd_addr_II[117]	(fmap_rd_addr_II[117]	),
    .\fmap_rd_addr_II[118]	(fmap_rd_addr_II[118]	),
    .\fmap_rd_addr_II[119]	(fmap_rd_addr_II[119]	),
    .\fmap_rd_addr_II[120]	(fmap_rd_addr_II[120]	),
    .\fmap_rd_addr_II[121]	(fmap_rd_addr_II[121]	),
    .\fmap_rd_addr_II[122]	(fmap_rd_addr_II[122]	),
    .\fmap_rd_addr_II[123]	(fmap_rd_addr_II[123]	),
    .\fmap_rd_addr_II[124]	(fmap_rd_addr_II[124]	),
    .\fmap_rd_addr_II[125]	(fmap_rd_addr_II[125]	),
    .\fmap_rd_addr_II[126]	(fmap_rd_addr_II[126]	),
    .\fmap_rd_addr_II[127]	(fmap_rd_addr_II[127]	),
    .\fmap_rd_addr_II[128]	(fmap_rd_addr_II[128]	),
    .\fmap_rd_addr_II[129]	(fmap_rd_addr_II[129]	),
    .\fmap_rd_addr_II[130]	(fmap_rd_addr_II[130]	),
    .\fmap_rd_addr_II[131]	(fmap_rd_addr_II[131]	),
    .\fmap_rd_addr_II[132]	(fmap_rd_addr_II[132]	),
    .\fmap_rd_addr_II[133]	(fmap_rd_addr_II[133]	),
    .\fmap_rd_addr_II[134]	(fmap_rd_addr_II[134]	),
    .\fmap_rd_addr_II[135]	(fmap_rd_addr_II[135]	),
    .\fmap_rd_addr_II[136]	(fmap_rd_addr_II[136]	),
    .\fmap_rd_addr_II[137]	(fmap_rd_addr_II[137]	),
    .\fmap_rd_addr_II[138]	(fmap_rd_addr_II[138]	),
    .\fmap_rd_addr_II[139]	(fmap_rd_addr_II[139]	),
    .\fmap_rd_addr_II[140]	(fmap_rd_addr_II[140]	),
    .\fmap_rd_addr_II[141]	(fmap_rd_addr_II[141]	),
    .\fmap_rd_addr_II[142]	(fmap_rd_addr_II[142]	),
    .\fmap_rd_addr_II[143]	(fmap_rd_addr_II[143]	),

    .\fmap_rd_addr_III[0]	(fmap_rd_addr_III[0]	),
    .\fmap_rd_addr_III[1]	(fmap_rd_addr_III[1]	),
    .\fmap_rd_addr_III[2]	(fmap_rd_addr_III[2]	),
    .\fmap_rd_addr_III[3]	(fmap_rd_addr_III[3]	),
    .\fmap_rd_addr_III[4]	(fmap_rd_addr_III[4]	),
    .\fmap_rd_addr_III[5]	(fmap_rd_addr_III[5]	),
    .\fmap_rd_addr_III[6]	(fmap_rd_addr_III[6]	),
    .\fmap_rd_addr_III[7]	(fmap_rd_addr_III[7]	),
    .\fmap_rd_addr_III[8]	(fmap_rd_addr_III[8]	),
    .\fmap_rd_addr_III[9]	(fmap_rd_addr_III[9]	),
    .\fmap_rd_addr_III[10]	(fmap_rd_addr_III[10]	),
    .\fmap_rd_addr_III[11]	(fmap_rd_addr_III[11]	),
    .\fmap_rd_addr_III[12]	(fmap_rd_addr_III[12]	),
    .\fmap_rd_addr_III[13]	(fmap_rd_addr_III[13]	),
    .\fmap_rd_addr_III[14]	(fmap_rd_addr_III[14]	),
    .\fmap_rd_addr_III[15]	(fmap_rd_addr_III[15]	),
    .\fmap_rd_addr_III[16]	(fmap_rd_addr_III[16]	),
    .\fmap_rd_addr_III[17]	(fmap_rd_addr_III[17]	),
    .\fmap_rd_addr_III[18]	(fmap_rd_addr_III[18]	),
    .\fmap_rd_addr_III[19]	(fmap_rd_addr_III[19]	),
    .\fmap_rd_addr_III[20]	(fmap_rd_addr_III[20]	),
    .\fmap_rd_addr_III[21]	(fmap_rd_addr_III[21]	),
    .\fmap_rd_addr_III[22]	(fmap_rd_addr_III[22]	),
    .\fmap_rd_addr_III[23]	(fmap_rd_addr_III[23]	),
    .\fmap_rd_addr_III[24]	(fmap_rd_addr_III[24]	),
    .\fmap_rd_addr_III[25]	(fmap_rd_addr_III[25]	),
    .\fmap_rd_addr_III[26]	(fmap_rd_addr_III[26]	),
    .\fmap_rd_addr_III[27]	(fmap_rd_addr_III[27]	),
    .\fmap_rd_addr_III[28]	(fmap_rd_addr_III[28]	),
    .\fmap_rd_addr_III[29]	(fmap_rd_addr_III[29]	),
    .\fmap_rd_addr_III[30]	(fmap_rd_addr_III[30]	),
    .\fmap_rd_addr_III[31]	(fmap_rd_addr_III[31]	),
    .\fmap_rd_addr_III[32]	(fmap_rd_addr_III[32]	),
    .\fmap_rd_addr_III[33]	(fmap_rd_addr_III[33]	),
    .\fmap_rd_addr_III[34]	(fmap_rd_addr_III[34]	),
    .\fmap_rd_addr_III[35]	(fmap_rd_addr_III[35]	),
    .\fmap_rd_addr_III[36]	(fmap_rd_addr_III[36]	),
    .\fmap_rd_addr_III[37]	(fmap_rd_addr_III[37]	),
    .\fmap_rd_addr_III[38]	(fmap_rd_addr_III[38]	),
    .\fmap_rd_addr_III[39]	(fmap_rd_addr_III[39]	),
    .\fmap_rd_addr_III[40]	(fmap_rd_addr_III[40]	),
    .\fmap_rd_addr_III[41]	(fmap_rd_addr_III[41]	),
    .\fmap_rd_addr_III[42]	(fmap_rd_addr_III[42]	),
    .\fmap_rd_addr_III[43]	(fmap_rd_addr_III[43]	),
    .\fmap_rd_addr_III[44]	(fmap_rd_addr_III[44]	),
    .\fmap_rd_addr_III[45]	(fmap_rd_addr_III[45]	),
    .\fmap_rd_addr_III[46]	(fmap_rd_addr_III[46]	),
    .\fmap_rd_addr_III[47]	(fmap_rd_addr_III[47]	),
    .\fmap_rd_addr_III[48]	(fmap_rd_addr_III[48]	),
    .\fmap_rd_addr_III[49]	(fmap_rd_addr_III[49]	),
    .\fmap_rd_addr_III[50]	(fmap_rd_addr_III[50]	),
    .\fmap_rd_addr_III[51]	(fmap_rd_addr_III[51]	),
    .\fmap_rd_addr_III[52]	(fmap_rd_addr_III[52]	),
    .\fmap_rd_addr_III[53]	(fmap_rd_addr_III[53]	),
    .\fmap_rd_addr_III[54]	(fmap_rd_addr_III[54]	),
    .\fmap_rd_addr_III[55]	(fmap_rd_addr_III[55]	),
    .\fmap_rd_addr_III[56]	(fmap_rd_addr_III[56]	),
    .\fmap_rd_addr_III[57]	(fmap_rd_addr_III[57]	),
    .\fmap_rd_addr_III[58]	(fmap_rd_addr_III[58]	),
    .\fmap_rd_addr_III[59]	(fmap_rd_addr_III[59]	),
    .\fmap_rd_addr_III[60]	(fmap_rd_addr_III[60]	),
    .\fmap_rd_addr_III[61]	(fmap_rd_addr_III[61]	),
    .\fmap_rd_addr_III[62]	(fmap_rd_addr_III[62]	),
    .\fmap_rd_addr_III[63]	(fmap_rd_addr_III[63]	),

    .\fmap_wr_addr_III[0]	(fmap_wr_addr_III[0]	),
    .\fmap_wr_addr_III[1]	(fmap_wr_addr_III[1]	),
    .\fmap_wr_addr_III[2]	(fmap_wr_addr_III[2]	),
    .\fmap_wr_addr_III[3]	(fmap_wr_addr_III[3]	),
    .\fmap_wr_addr_III[4]	(fmap_wr_addr_III[4]	),
    .\fmap_wr_addr_III[5]	(fmap_wr_addr_III[5]	),
    .\fmap_wr_addr_III[6]	(fmap_wr_addr_III[6]	),
    .\fmap_wr_addr_III[7]	(fmap_wr_addr_III[7]	),
    .\fmap_wr_addr_III[8]	(fmap_wr_addr_III[8]	),
    .\fmap_wr_addr_III[9]	(fmap_wr_addr_III[9]	),
    .\fmap_wr_addr_III[10]	(fmap_wr_addr_III[10]	),
    .\fmap_wr_addr_III[11]	(fmap_wr_addr_III[11]	),
    .\fmap_wr_addr_III[12]	(fmap_wr_addr_III[12]	),
    .\fmap_wr_addr_III[13]	(fmap_wr_addr_III[13]	),
    .\fmap_wr_addr_III[14]	(fmap_wr_addr_III[14]	),
    .\fmap_wr_addr_III[15]	(fmap_wr_addr_III[15]	),
    .\fmap_wr_addr_III[16]	(fmap_wr_addr_III[16]	),
    .\fmap_wr_addr_III[17]	(fmap_wr_addr_III[17]	),
    .\fmap_wr_addr_III[18]	(fmap_wr_addr_III[18]	),
    .\fmap_wr_addr_III[19]	(fmap_wr_addr_III[19]	),
    .\fmap_wr_addr_III[20]	(fmap_wr_addr_III[20]	),
    .\fmap_wr_addr_III[21]	(fmap_wr_addr_III[21]	),
    .\fmap_wr_addr_III[22]	(fmap_wr_addr_III[22]	),
    .\fmap_wr_addr_III[23]	(fmap_wr_addr_III[23]	),
    .\fmap_wr_addr_III[24]	(fmap_wr_addr_III[24]	),
    .\fmap_wr_addr_III[25]	(fmap_wr_addr_III[25]	),
    .\fmap_wr_addr_III[26]	(fmap_wr_addr_III[26]	),
    .\fmap_wr_addr_III[27]	(fmap_wr_addr_III[27]	),
    .\fmap_wr_addr_III[28]	(fmap_wr_addr_III[28]	),
    .\fmap_wr_addr_III[29]	(fmap_wr_addr_III[29]	),
    .\fmap_wr_addr_III[30]	(fmap_wr_addr_III[30]	),
    .\fmap_wr_addr_III[31]	(fmap_wr_addr_III[31]	),
    .\fmap_wr_addr_III[32]	(fmap_wr_addr_III[32]	),
    .\fmap_wr_addr_III[33]	(fmap_wr_addr_III[33]	),
    .\fmap_wr_addr_III[34]	(fmap_wr_addr_III[34]	),
    .\fmap_wr_addr_III[35]	(fmap_wr_addr_III[35]	),
    .\fmap_wr_addr_III[36]	(fmap_wr_addr_III[36]	),
    .\fmap_wr_addr_III[37]	(fmap_wr_addr_III[37]	),
    .\fmap_wr_addr_III[38]	(fmap_wr_addr_III[38]	),
    .\fmap_wr_addr_III[39]	(fmap_wr_addr_III[39]	),
    .\fmap_wr_addr_III[40]	(fmap_wr_addr_III[40]	),
    .\fmap_wr_addr_III[41]	(fmap_wr_addr_III[41]	),
    .\fmap_wr_addr_III[42]	(fmap_wr_addr_III[42]	),
    .\fmap_wr_addr_III[43]	(fmap_wr_addr_III[43]	),
    .\fmap_wr_addr_III[44]	(fmap_wr_addr_III[44]	),
    .\fmap_wr_addr_III[45]	(fmap_wr_addr_III[45]	),
    .\fmap_wr_addr_III[46]	(fmap_wr_addr_III[46]	),
    .\fmap_wr_addr_III[47]	(fmap_wr_addr_III[47]	),
    .\fmap_wr_addr_III[48]	(fmap_wr_addr_III[48]	),
    .\fmap_wr_addr_III[49]	(fmap_wr_addr_III[49]	),
    .\fmap_wr_addr_III[50]	(fmap_wr_addr_III[50]	),
    .\fmap_wr_addr_III[51]	(fmap_wr_addr_III[51]	),
    .\fmap_wr_addr_III[52]	(fmap_wr_addr_III[52]	),
    .\fmap_wr_addr_III[53]	(fmap_wr_addr_III[53]	),
    .\fmap_wr_addr_III[54]	(fmap_wr_addr_III[54]	),
    .\fmap_wr_addr_III[55]	(fmap_wr_addr_III[55]	),
    .\fmap_wr_addr_III[56]	(fmap_wr_addr_III[56]	),
    .\fmap_wr_addr_III[57]	(fmap_wr_addr_III[57]	),
    .\fmap_wr_addr_III[58]	(fmap_wr_addr_III[58]	),
    .\fmap_wr_addr_III[59]	(fmap_wr_addr_III[59]	),
    .\fmap_wr_addr_III[60]	(fmap_wr_addr_III[60]	),
    .\fmap_wr_addr_III[61]	(fmap_wr_addr_III[61]	),
    .\fmap_wr_addr_III[62]	(fmap_wr_addr_III[62]	),
    .\fmap_wr_addr_III[63]	(fmap_wr_addr_III[63]	),

    .\fmap_wr_en_III[0]	(fmap_wr_en_III[0]	),
    .\fmap_wr_en_III[1]	(fmap_wr_en_III[1]	),
    .\fmap_wr_en_III[2]	(fmap_wr_en_III[2]	),
    .\fmap_wr_en_III[3]	(fmap_wr_en_III[3]	),
    .\fmap_wr_en_III[4]	(fmap_wr_en_III[4]	),
    .\fmap_wr_en_III[5]	(fmap_wr_en_III[5]	),
    .\fmap_wr_en_III[6]	(fmap_wr_en_III[6]	),
    .\fmap_wr_en_III[7]	(fmap_wr_en_III[7]	),
    .\fmap_wr_en_III[8]	(fmap_wr_en_III[8]	),
    .\fmap_wr_en_III[9]	(fmap_wr_en_III[9]	),
    .\fmap_wr_en_III[10]	(fmap_wr_en_III[10]	),
    .\fmap_wr_en_III[11]	(fmap_wr_en_III[11]	),
    .\fmap_wr_en_III[12]	(fmap_wr_en_III[12]	),
    .\fmap_wr_en_III[13]	(fmap_wr_en_III[13]	),
    .\fmap_wr_en_III[14]	(fmap_wr_en_III[14]	),
    .\fmap_wr_en_III[15]	(fmap_wr_en_III[15]	),
    .\fmap_wr_en_III[16]	(fmap_wr_en_III[16]	),
    .\fmap_wr_en_III[17]	(fmap_wr_en_III[17]	),
    .\fmap_wr_en_III[18]	(fmap_wr_en_III[18]	),
    .\fmap_wr_en_III[19]	(fmap_wr_en_III[19]	),
    .\fmap_wr_en_III[20]	(fmap_wr_en_III[20]	),
    .\fmap_wr_en_III[21]	(fmap_wr_en_III[21]	),
    .\fmap_wr_en_III[22]	(fmap_wr_en_III[22]	),
    .\fmap_wr_en_III[23]	(fmap_wr_en_III[23]	),
    .\fmap_wr_en_III[24]	(fmap_wr_en_III[24]	),
    .\fmap_wr_en_III[25]	(fmap_wr_en_III[25]	),
    .\fmap_wr_en_III[26]	(fmap_wr_en_III[26]	),
    .\fmap_wr_en_III[27]	(fmap_wr_en_III[27]	),
    .\fmap_wr_en_III[28]	(fmap_wr_en_III[28]	),
    .\fmap_wr_en_III[29]	(fmap_wr_en_III[29]	),
    .\fmap_wr_en_III[30]	(fmap_wr_en_III[30]	),
    .\fmap_wr_en_III[31]	(fmap_wr_en_III[31]	),
    .\fmap_wr_en_III[32]	(fmap_wr_en_III[32]	),
    .\fmap_wr_en_III[33]	(fmap_wr_en_III[33]	),
    .\fmap_wr_en_III[34]	(fmap_wr_en_III[34]	),
    .\fmap_wr_en_III[35]	(fmap_wr_en_III[35]	),
    .\fmap_wr_en_III[36]	(fmap_wr_en_III[36]	),
    .\fmap_wr_en_III[37]	(fmap_wr_en_III[37]	),
    .\fmap_wr_en_III[38]	(fmap_wr_en_III[38]	),
    .\fmap_wr_en_III[39]	(fmap_wr_en_III[39]	),
    .\fmap_wr_en_III[40]	(fmap_wr_en_III[40]	),
    .\fmap_wr_en_III[41]	(fmap_wr_en_III[41]	),
    .\fmap_wr_en_III[42]	(fmap_wr_en_III[42]	),
    .\fmap_wr_en_III[43]	(fmap_wr_en_III[43]	),
    .\fmap_wr_en_III[44]	(fmap_wr_en_III[44]	),
    .\fmap_wr_en_III[45]	(fmap_wr_en_III[45]	),
    .\fmap_wr_en_III[46]	(fmap_wr_en_III[46]	),
    .\fmap_wr_en_III[47]	(fmap_wr_en_III[47]	),
    .\fmap_wr_en_III[48]	(fmap_wr_en_III[48]	),
    .\fmap_wr_en_III[49]	(fmap_wr_en_III[49]	),
    .\fmap_wr_en_III[50]	(fmap_wr_en_III[50]	),
    .\fmap_wr_en_III[51]	(fmap_wr_en_III[51]	),
    .\fmap_wr_en_III[52]	(fmap_wr_en_III[52]	),
    .\fmap_wr_en_III[53]	(fmap_wr_en_III[53]	),
    .\fmap_wr_en_III[54]	(fmap_wr_en_III[54]	),
    .\fmap_wr_en_III[55]	(fmap_wr_en_III[55]	),
    .\fmap_wr_en_III[56]	(fmap_wr_en_III[56]	),
    .\fmap_wr_en_III[57]	(fmap_wr_en_III[57]	),
    .\fmap_wr_en_III[58]	(fmap_wr_en_III[58]	),
    .\fmap_wr_en_III[59]	(fmap_wr_en_III[59]	),
    .\fmap_wr_en_III[60]	(fmap_wr_en_III[60]	),
    .\fmap_wr_en_III[61]	(fmap_wr_en_III[61]	),
    .\fmap_wr_en_III[62]	(fmap_wr_en_III[62]	),
    .\fmap_wr_en_III[63]	(fmap_wr_en_III[63]	),

    .\fmap_wr_data_III[0]	(fmap_wr_data_III[0]	),
    .\fmap_wr_data_III[1]	(fmap_wr_data_III[1]	),
    .\fmap_wr_data_III[2]	(fmap_wr_data_III[2]	),
    .\fmap_wr_data_III[3]	(fmap_wr_data_III[3]	),
    .\fmap_wr_data_III[4]	(fmap_wr_data_III[4]	),
    .\fmap_wr_data_III[5]	(fmap_wr_data_III[5]	),
    .\fmap_wr_data_III[6]	(fmap_wr_data_III[6]	),
    .\fmap_wr_data_III[7]	(fmap_wr_data_III[7]	),
    .\fmap_wr_data_III[8]	(fmap_wr_data_III[8]	),
    .\fmap_wr_data_III[9]	(fmap_wr_data_III[9]	),
    .\fmap_wr_data_III[10]	(fmap_wr_data_III[10]	),
    .\fmap_wr_data_III[11]	(fmap_wr_data_III[11]	),
    .\fmap_wr_data_III[12]	(fmap_wr_data_III[12]	),
    .\fmap_wr_data_III[13]	(fmap_wr_data_III[13]	),
    .\fmap_wr_data_III[14]	(fmap_wr_data_III[14]	),
    .\fmap_wr_data_III[15]	(fmap_wr_data_III[15]	),
    .\fmap_wr_data_III[16]	(fmap_wr_data_III[16]	),
    .\fmap_wr_data_III[17]	(fmap_wr_data_III[17]	),
    .\fmap_wr_data_III[18]	(fmap_wr_data_III[18]	),
    .\fmap_wr_data_III[19]	(fmap_wr_data_III[19]	),
    .\fmap_wr_data_III[20]	(fmap_wr_data_III[20]	),
    .\fmap_wr_data_III[21]	(fmap_wr_data_III[21]	),
    .\fmap_wr_data_III[22]	(fmap_wr_data_III[22]	),
    .\fmap_wr_data_III[23]	(fmap_wr_data_III[23]	),
    .\fmap_wr_data_III[24]	(fmap_wr_data_III[24]	),
    .\fmap_wr_data_III[25]	(fmap_wr_data_III[25]	),
    .\fmap_wr_data_III[26]	(fmap_wr_data_III[26]	),
    .\fmap_wr_data_III[27]	(fmap_wr_data_III[27]	),
    .\fmap_wr_data_III[28]	(fmap_wr_data_III[28]	),
    .\fmap_wr_data_III[29]	(fmap_wr_data_III[29]	),
    .\fmap_wr_data_III[30]	(fmap_wr_data_III[30]	),
    .\fmap_wr_data_III[31]	(fmap_wr_data_III[31]	),
    .\fmap_wr_data_III[32]	(fmap_wr_data_III[32]	),
    .\fmap_wr_data_III[33]	(fmap_wr_data_III[33]	),
    .\fmap_wr_data_III[34]	(fmap_wr_data_III[34]	),
    .\fmap_wr_data_III[35]	(fmap_wr_data_III[35]	),
    .\fmap_wr_data_III[36]	(fmap_wr_data_III[36]	),
    .\fmap_wr_data_III[37]	(fmap_wr_data_III[37]	),
    .\fmap_wr_data_III[38]	(fmap_wr_data_III[38]	),
    .\fmap_wr_data_III[39]	(fmap_wr_data_III[39]	),
    .\fmap_wr_data_III[40]	(fmap_wr_data_III[40]	),
    .\fmap_wr_data_III[41]	(fmap_wr_data_III[41]	),
    .\fmap_wr_data_III[42]	(fmap_wr_data_III[42]	),
    .\fmap_wr_data_III[43]	(fmap_wr_data_III[43]	),
    .\fmap_wr_data_III[44]	(fmap_wr_data_III[44]	),
    .\fmap_wr_data_III[45]	(fmap_wr_data_III[45]	),
    .\fmap_wr_data_III[46]	(fmap_wr_data_III[46]	),
    .\fmap_wr_data_III[47]	(fmap_wr_data_III[47]	),
    .\fmap_wr_data_III[48]	(fmap_wr_data_III[48]	),
    .\fmap_wr_data_III[49]	(fmap_wr_data_III[49]	),
    .\fmap_wr_data_III[50]	(fmap_wr_data_III[50]	),
    .\fmap_wr_data_III[51]	(fmap_wr_data_III[51]	),
    .\fmap_wr_data_III[52]	(fmap_wr_data_III[52]	),
    .\fmap_wr_data_III[53]	(fmap_wr_data_III[53]	),
    .\fmap_wr_data_III[54]	(fmap_wr_data_III[54]	),
    .\fmap_wr_data_III[55]	(fmap_wr_data_III[55]	),
    .\fmap_wr_data_III[56]	(fmap_wr_data_III[56]	),
    .\fmap_wr_data_III[57]	(fmap_wr_data_III[57]	),
    .\fmap_wr_data_III[58]	(fmap_wr_data_III[58]	),
    .\fmap_wr_data_III[59]	(fmap_wr_data_III[59]	),
    .\fmap_wr_data_III[60]	(fmap_wr_data_III[60]	),
    .\fmap_wr_data_III[61]	(fmap_wr_data_III[61]	),
    .\fmap_wr_data_III[62]	(fmap_wr_data_III[62]	),
    .\fmap_wr_data_III[63]	(fmap_wr_data_III[63]	),

    .\fmap_rd_data_III[0]	(fmap_rd_data_III[0]	),
    .\fmap_rd_data_III[1]	(fmap_rd_data_III[1]	),
    .\fmap_rd_data_III[2]	(fmap_rd_data_III[2]	),
    .\fmap_rd_data_III[3]	(fmap_rd_data_III[3]	),
    .\fmap_rd_data_III[4]	(fmap_rd_data_III[4]	),
    .\fmap_rd_data_III[5]	(fmap_rd_data_III[5]	),
    .\fmap_rd_data_III[6]	(fmap_rd_data_III[6]	),
    .\fmap_rd_data_III[7]	(fmap_rd_data_III[7]	),
    .\fmap_rd_data_III[8]	(fmap_rd_data_III[8]	),
    .\fmap_rd_data_III[9]	(fmap_rd_data_III[9]	),
    .\fmap_rd_data_III[10]	(fmap_rd_data_III[10]	),
    .\fmap_rd_data_III[11]	(fmap_rd_data_III[11]	),
    .\fmap_rd_data_III[12]	(fmap_rd_data_III[12]	),
    .\fmap_rd_data_III[13]	(fmap_rd_data_III[13]	),
    .\fmap_rd_data_III[14]	(fmap_rd_data_III[14]	),
    .\fmap_rd_data_III[15]	(fmap_rd_data_III[15]	),
    .\fmap_rd_data_III[16]	(fmap_rd_data_III[16]	),
    .\fmap_rd_data_III[17]	(fmap_rd_data_III[17]	),
    .\fmap_rd_data_III[18]	(fmap_rd_data_III[18]	),
    .\fmap_rd_data_III[19]	(fmap_rd_data_III[19]	),
    .\fmap_rd_data_III[20]	(fmap_rd_data_III[20]	),
    .\fmap_rd_data_III[21]	(fmap_rd_data_III[21]	),
    .\fmap_rd_data_III[22]	(fmap_rd_data_III[22]	),
    .\fmap_rd_data_III[23]	(fmap_rd_data_III[23]	),
    .\fmap_rd_data_III[24]	(fmap_rd_data_III[24]	),
    .\fmap_rd_data_III[25]	(fmap_rd_data_III[25]	),
    .\fmap_rd_data_III[26]	(fmap_rd_data_III[26]	),
    .\fmap_rd_data_III[27]	(fmap_rd_data_III[27]	),
    .\fmap_rd_data_III[28]	(fmap_rd_data_III[28]	),
    .\fmap_rd_data_III[29]	(fmap_rd_data_III[29]	),
    .\fmap_rd_data_III[30]	(fmap_rd_data_III[30]	),
    .\fmap_rd_data_III[31]	(fmap_rd_data_III[31]	),
    .\fmap_rd_data_III[32]	(fmap_rd_data_III[32]	),
    .\fmap_rd_data_III[33]	(fmap_rd_data_III[33]	),
    .\fmap_rd_data_III[34]	(fmap_rd_data_III[34]	),
    .\fmap_rd_data_III[35]	(fmap_rd_data_III[35]	),
    .\fmap_rd_data_III[36]	(fmap_rd_data_III[36]	),
    .\fmap_rd_data_III[37]	(fmap_rd_data_III[37]	),
    .\fmap_rd_data_III[38]	(fmap_rd_data_III[38]	),
    .\fmap_rd_data_III[39]	(fmap_rd_data_III[39]	),
    .\fmap_rd_data_III[40]	(fmap_rd_data_III[40]	),
    .\fmap_rd_data_III[41]	(fmap_rd_data_III[41]	),
    .\fmap_rd_data_III[42]	(fmap_rd_data_III[42]	),
    .\fmap_rd_data_III[43]	(fmap_rd_data_III[43]	),
    .\fmap_rd_data_III[44]	(fmap_rd_data_III[44]	),
    .\fmap_rd_data_III[45]	(fmap_rd_data_III[45]	),
    .\fmap_rd_data_III[46]	(fmap_rd_data_III[46]	),
    .\fmap_rd_data_III[47]	(fmap_rd_data_III[47]	),
    .\fmap_rd_data_III[48]	(fmap_rd_data_III[48]	),
    .\fmap_rd_data_III[49]	(fmap_rd_data_III[49]	),
    .\fmap_rd_data_III[50]	(fmap_rd_data_III[50]	),
    .\fmap_rd_data_III[51]	(fmap_rd_data_III[51]	),
    .\fmap_rd_data_III[52]	(fmap_rd_data_III[52]	),
    .\fmap_rd_data_III[53]	(fmap_rd_data_III[53]	),
    .\fmap_rd_data_III[54]	(fmap_rd_data_III[54]	),
    .\fmap_rd_data_III[55]	(fmap_rd_data_III[55]	),
    .\fmap_rd_data_III[56]	(fmap_rd_data_III[56]	),
    .\fmap_rd_data_III[57]	(fmap_rd_data_III[57]	),
    .\fmap_rd_data_III[58]	(fmap_rd_data_III[58]	),
    .\fmap_rd_data_III[59]	(fmap_rd_data_III[59]	),
    .\fmap_rd_data_III[60]	(fmap_rd_data_III[60]	),
    .\fmap_rd_data_III[61]	(fmap_rd_data_III[61]	),
    .\fmap_rd_data_III[62]	(fmap_rd_data_III[62]	),
    .\fmap_rd_data_III[63]	(fmap_rd_data_III[63]	),

    // Classification. (fmap III -> FC7 -> 10 registers -> apply max -> get "digit_o" right here)
    .digit_o       (digit_o),
    .digit_o_valid (digit_o_valid)
    
);

// Line buffer memory
ff_line_buffer_groups #(
    .LINE_BUF_GROUPS(LINE_BUF_GROUPS),
    .LINE_BUFS_PER_GROUP(LINE_BUFS_PER_GROUP),
    .LINE_BUF_ADDR_BITS(LINE_BUF_ADDR_BITS),
    .D_WIDTH(D_WIDTH),
    .LINE_BUF_DEPTH(LINE_BUF_DEPTH)
)
ff_line_buffer_groups_u 
(
    .clk(clk),
    .line_buffer_rd_addr(line_buffer_rd_addr),
    .line_buffer_wr_addr(line_buffer_wr_addr),
    .line_buffer_wr_data(line_buffer_wr_data),
    .line_buffer_wr_en(line_buffer_wr_en),
    .line_buffer_rd_data(line_buffer_rd_data)  
);

// Fmap memory
fmap_I #(
    .ADDR_WIDTH(FMAP_I_ADDR_BITS),
    .DATA_WIDTH(D_WIDTH),
    .DEPTH(FMAP_I_DEPTH)
)
fmap_I_u 
(
    .clk(clk),
    .wr_addr_1(fmap_wr_addr_I[0]),
    .wr_addr_2(fmap_wr_addr_I[1]),
    .wr_addr_3(fmap_wr_addr_I[2]),
    .wr_addr_4(fmap_wr_addr_I[3]),
    .wr_addr_5(fmap_wr_addr_I[4]),
    .wr_addr_6(fmap_wr_addr_I[5]),
    .wr_addr_7(fmap_wr_addr_I[6]),
    .wr_addr_8(fmap_wr_addr_I[7]),
    .wr_addr_9(fmap_wr_addr_I[8]),
    .wr_addr_10(fmap_wr_addr_I[9]),
    .wr_addr_11(fmap_wr_addr_I[10]),
    .wr_addr_12(fmap_wr_addr_I[11]),
    .wr_addr_13(fmap_wr_addr_I[12]),
    .wr_addr_14(fmap_wr_addr_I[13]),
    .wr_addr_15(fmap_wr_addr_I[14]),
    .wr_addr_16(fmap_wr_addr_I[15]),
    .rd_addr_1(fmap_rd_addr_I[0]),
    .rd_addr_2(fmap_rd_addr_I[1]),
    .rd_addr_3(fmap_rd_addr_I[2]),
    .rd_addr_4(fmap_rd_addr_I[3]),
    .rd_addr_5(fmap_rd_addr_I[4]),
    .rd_addr_6(fmap_rd_addr_I[5]),
    .rd_addr_7(fmap_rd_addr_I[6]),
    .rd_addr_8(fmap_rd_addr_I[7]),
    .rd_addr_9(fmap_rd_addr_I[8]),
    .rd_addr_10(fmap_rd_addr_I[9]),
    .rd_addr_11(fmap_rd_addr_I[10]),
    .rd_addr_12(fmap_rd_addr_I[11]),
    .rd_addr_13(fmap_rd_addr_I[12]),
    .rd_addr_14(fmap_rd_addr_I[13]),
    .rd_addr_15(fmap_rd_addr_I[14]),
    .rd_addr_16(fmap_rd_addr_I[15]),
    .wr_en_1(fmap_wr_en_I[0]),
    .wr_en_2(fmap_wr_en_I[1]),
    .wr_en_3(fmap_wr_en_I[2]),
    .wr_en_4(fmap_wr_en_I[3]),
    .wr_en_5(fmap_wr_en_I[4]),
    .wr_en_6(fmap_wr_en_I[5]),
    .wr_en_7(fmap_wr_en_I[6]),
    .wr_en_8(fmap_wr_en_I[7]),
    .wr_en_9(fmap_wr_en_I[8]),
    .wr_en_10(fmap_wr_en_I[9]),
    .wr_en_11(fmap_wr_en_I[10]),
    .wr_en_12(fmap_wr_en_I[11]),
    .wr_en_13(fmap_wr_en_I[12]),
    .wr_en_14(fmap_wr_en_I[13]),
    .wr_en_15(fmap_wr_en_I[14]),
    .wr_en_16(fmap_wr_en_I[15]),
    .wr_data_1(fmap_wr_data_I[0]),
    .wr_data_2(fmap_wr_data_I[1]),
    .wr_data_3(fmap_wr_data_I[2]),
    .wr_data_4(fmap_wr_data_I[3]),
    .wr_data_5(fmap_wr_data_I[4]),
    .wr_data_6(fmap_wr_data_I[5]),
    .wr_data_7(fmap_wr_data_I[6]),
    .wr_data_8(fmap_wr_data_I[7]),
    .wr_data_9(fmap_wr_data_I[8]),
    .wr_data_10(fmap_wr_data_I[9]),
    .wr_data_11(fmap_wr_data_I[10]),
    .wr_data_12(fmap_wr_data_I[11]),
    .wr_data_13(fmap_wr_data_I[12]),
    .wr_data_14(fmap_wr_data_I[13]),
    .wr_data_15(fmap_wr_data_I[14]),
    .wr_data_16(fmap_wr_data_I[15]),
    .rd_data_1(fmap_rd_data_I[0]),
    .rd_data_2(fmap_rd_data_I[1]),
    .rd_data_3(fmap_rd_data_I[2]),
    .rd_data_4(fmap_rd_data_I[3]),
    .rd_data_5(fmap_rd_data_I[4]),
    .rd_data_6(fmap_rd_data_I[5]),
    .rd_data_7(fmap_rd_data_I[6]),
    .rd_data_8(fmap_rd_data_I[7]),
    .rd_data_9(fmap_rd_data_I[8]),
    .rd_data_10(fmap_rd_data_I[9]),
    .rd_data_11(fmap_rd_data_I[10]),
    .rd_data_12(fmap_rd_data_I[11]),
    .rd_data_13(fmap_rd_data_I[12]),
    .rd_data_14(fmap_rd_data_I[13]),
    .rd_data_15(fmap_rd_data_I[14]),
    .rd_data_16(fmap_rd_data_I[15])
);

fmap_II fmap_II_u 
(
    .clk(clk),
    .fmap_wr_addr(fmap_wr_addr_II),
    .fmap_rd_addr(fmap_rd_addr_II),
    .fmap_wr_en(fmap_wr_en_II),
    .fmap_wr_data(fmap_wr_data_II),
    .fmap_rd_data(fmap_rd_data_II)
);

fmap_III fmap_III_u 
(
    .clk(clk),
    .fmap_wr_addr(fmap_wr_addr_III),
    .fmap_rd_addr(fmap_rd_addr_III),
    .fmap_wr_en(fmap_wr_en_III),
    .fmap_wr_data(fmap_wr_data_III),
    .fmap_rd_data(fmap_rd_data_III)
);

// Bias memory
bi_mem0 bi_mem0_u 
(
    .clk(clk),
    .addr_a(bi_addr_a),
    .addr_b(bi_addr_b),
    .q_a(bi_q_a),
    .q_b(bi_q_b)
);

// Weights memory
wt_mem0 wt_mem0_u (
    .clk(clk),
    .addr_a(addr_a[0]),
    .addr_b(addr_b[0]),
    .q_a(q_a[0]),
    .q_b(q_b[0])
);

wt_mem1 wt_mem1_u (
    .clk(clk),
    .addr_a(addr_a[1]),
    .addr_b(addr_b[1]),
    .q_a(q_a[1]),
    .q_b(q_b[1])
);

wt_mem2 wt_mem2_u (
    .clk(clk),
    .addr_a(addr_a[2]),
    .addr_b(addr_b[2]),
    .q_a(q_a[2]),
    .q_b(q_b[2])
);

wt_mem3 wt_mem3_u (
    .clk(clk),
    .addr_a(addr_a[3]),
    .addr_b(addr_b[3]),
    .q_a(q_a[3]),
    .q_b(q_b[3])
);

wt_mem4 wt_mem4_u (
    .clk(clk),
    .addr_a(addr_a[4]),
    .addr_b(addr_b[4]),
    .q_a(q_a[4]),
    .q_b(q_b[4])
);

wt_mem5 wt_mem5_u (
    .clk(clk),
    .addr_a(addr_a[5]),
    .addr_b(addr_b[5]),
    .q_a(q_a[5]),
    .q_b(q_b[5])
);

wt_mem6 wt_mem6_u (
    .clk(clk),
    .addr_a(addr_a[6]),
    .addr_b(addr_b[6]),
    .q_a(q_a[6]),
    .q_b(q_b[6])
);

wt_mem7 wt_mem7_u (
    .clk(clk),
    .addr_a(addr_a[7]),
    .addr_b(addr_b[7]),
    .q_a(q_a[7]),
    .q_b(q_b[7])
);


endmodule
