`timescale 1ns/1ns

module wt_mem0 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h10a71653eefa15980348fe98e491e22819d6;
mem[1] = 144'h1346f6e1082eee57ec73fe661a0aefb8f687;
mem[2] = 144'hf9a0e7e2fab4e4cfebbee32cef53ef4819c0;
mem[3] = 144'hee71fbe1fb88eaecf3e9ebd3ee921b1819e9;
mem[4] = 144'h134beef6ff2d0473184cea8aeb74e1ce1e46;
mem[5] = 144'he2100ad1fd7d03e2ec311ed4185ff79fea05;
mem[6] = 144'h07f50aa90c751c8ef24ee459eecf0ac5f045;
mem[7] = 144'hf456093002dae796fe9a09681c2608e302c9;
mem[8] = 144'h11111f170540eaa100c9e9a617071886ecbe;
mem[9] = 144'he7dfec18f208ed21e2b50274e95a08a30c7c;
mem[10] = 144'heb660167ed5ff704f57f19efe3a1eb3f0b3d;
mem[11] = 144'h18fee34913181322e4aa1c5a0effe5aa0bc2;
mem[12] = 144'he3cd0c92e5daf436e805e0431174e854fb0e;
mem[13] = 144'h1be310e40f99fd4e1099e6c7ef640f670b9f;
mem[14] = 144'he1e90e5a0eb8fafbf7c4047deb7115f5eb68;
mem[15] = 144'hfa59055800be068d034ce5450fff05550e0a;
mem[16] = 144'hf5d40f1ff9c61b9a093c0fa0e86a15111514;
mem[17] = 144'hf53ae7c91b85e9c01898f985f664e609e301;
mem[18] = 144'h0ab8e43d1b67eccdf99d144509350a70ffc3;
mem[19] = 144'he564f339e5f5ea7be085e936f4b702740861;
mem[20] = 144'h0aed04a206690008e7d4e38dedc60aaae390;
mem[21] = 144'he4beee20e91ff935e015f128e038ec1ceb32;
mem[22] = 144'h088ff2ad10fe02f0000404ddfc0010540f7f;
mem[23] = 144'hf1e71d4ceb0b0fd107b5e5c8ef2b066bf056;
mem[24] = 144'hf6d617aa1e820189f452e48e0d1108c90553;
mem[25] = 144'hecaf1859eb78ec7cfe271dfcf4ecf9d7fa09;
mem[26] = 144'hf3ae1d4ee0631257e71405ba2020ef10e6a7;
mem[27] = 144'h0f6414fc017c0c28f2bef4d814a4f3d51542;
mem[28] = 144'he29ff5340bbded36ee6b1d6ff93a1bbefbf3;
mem[29] = 144'h1318ef241e431f300cea1e29ea2df8030929;
mem[30] = 144'he75a03421796fd841352e308fcc10cbfedd0;
mem[31] = 144'h04b40cdafc9204af1307fdd1f260fc50f1df;
mem[32] = 144'h09e90a82e1a901f6e8781e95f5a6ea851f36;
mem[33] = 144'h133e005804e51ac1f9f906dae8ceeb35edc8;
mem[34] = 144'h1643fad6f05703bdf6f01b9019abff59fdfd;
mem[35] = 144'h1b4317010080f319f5ca16d4f5a3e8d7f898;
mem[36] = 144'hef90e5cf159609681e6615cd15ede158e340;
mem[37] = 144'h119fe3d1116606e7f131fe5d1cae1f220b86;
mem[38] = 144'hfc57f8d9111d0d4400cfe368f51a18bff104;
mem[39] = 144'h1e090537ffb2edc4f9b109aa10a3008e0f8b;
mem[40] = 144'h1d1d001c16101ea7172213e3e1f9ef2d07d8;
mem[41] = 144'heff1e32d0fd5f0320bd71e94111b077ef88f;
mem[42] = 144'hfe741c14ed2af778077dfc060a04f206e199;
mem[43] = 144'hf547eadcf0180ff01cf30507093f02c51a97;
mem[44] = 144'hff27068ee8ccf4ee03cdf616eb4a1007e933;
mem[45] = 144'hf31c000b049cffc5f1a7fa5b18f50230e0f4;
mem[46] = 144'h1200f3a1e384fd601d4d0eb0145df0f61410;
mem[47] = 144'h1451e556f4441ec8f5961ee41724ef1502eb;
mem[48] = 144'h1c25eea514f9feefe65811c80231e322ec33;
mem[49] = 144'hed0e09a3f5ad1f93edbcec88e5fdef85003b;
mem[50] = 144'h1ace0fcfe2c4063af84efe390cd4efc60935;
mem[51] = 144'h1b33e83aec97e53df034e7cbfeec189302cb;
mem[52] = 144'h089f0f77e9ab09d91517f8190b27008c1420;
mem[53] = 144'h03cc1187ea4cfdbb09d9fb9cfb870a16003f;
mem[54] = 144'heea9e97ee10aeb74ecca1d20ea9a1d1be173;
mem[55] = 144'h01751f9eff67f97206b0fc0ffeac1c7e117d;
mem[56] = 144'h040f1294e0c5f800e940eba3ed98ff4dfee1;
mem[57] = 144'he7adf065ed5804981f590a9d1cc1f6631e4b;
mem[58] = 144'hfc3fede5f5d9fcf4184110e01c4de0d8f58a;
mem[59] = 144'h1ef807f716571eb40e9bec27f002ffe1e7e4;
mem[60] = 144'hefd7e104efd5e1c4072109020cb7f9f9f453;
mem[61] = 144'hefb7f794feccec66e07ff3bee5ce068d0f9f;
mem[62] = 144'h18d5f4bd19acff6703270b4c1399f8e2152f;
mem[63] = 144'h1218e48be3f90213080de84cf037e195fcd7;
mem[64] = 144'he266ff25068ef9c018e3e24beffdf258ea85;
mem[65] = 144'h0184098e0872099e10d1f1cff8a504d815c0;
mem[66] = 144'he997ee39e37bf706f4330a381846fc001a9f;
mem[67] = 144'h17c80325f82dfd770022e51d0466f06bfb6c;
mem[68] = 144'h0ccb0e5cec01f247eb281b55f364fdde0a21;
mem[69] = 144'h03681cd61dc9ff84090412f3e19b12ec12fe;
mem[70] = 144'h01530a5ff87ce80ee33be5f6eea711dffe9f;
mem[71] = 144'he498e0c818da081eee1d1fd50ee1eebbf185;
mem[72] = 144'h02411dcafacffc251e76f6d1f7ca07851714;
mem[73] = 144'h1ef2050be6c1ef20ef2e19f6f2d0f8600648;
mem[74] = 144'h118aedd70db4fc7c1609e022e889e47319aa;
mem[75] = 144'he3241c5a0c5b1d90f8241e0715ee1244ee6e;
mem[76] = 144'hf896f0b41674ea81fc8d133d0353f6dd0aaa;
mem[77] = 144'hed48e168f606eeee1b6bff6bfc67e0081afe;
mem[78] = 144'heac6eaee0668fac717fcede2ef511fb1ff18;
mem[79] = 144'h01d60f85e9ea0fbc0ba5ea701cc608f6e981;
mem[80] = 144'h1acffa8c0fa0fb861f68128af1ae1c0c0be8;
mem[81] = 144'hf26c071918e8e050e973fa5ef904f4adebbe;
mem[82] = 144'h0c95e55af0a4e7fe1f9e065e03b4f489075d;
mem[83] = 144'he9221835012711c30f240f10ec63e37709e8;
mem[84] = 144'hf683fa07eaf507dc1cd7e611114a1539eb55;
mem[85] = 144'h1eed1d67f1fff59819e51e230b041ccbe197;
mem[86] = 144'h116e0165e4510b09f20aece50d4cf6570d7a;
mem[87] = 144'he105f3fa1ab402cf1ad20708e1e1e8fa1a6a;
mem[88] = 144'hf971fa52e788f588e1dbe7c3e13b02ec1632;
mem[89] = 144'h0209f62fefc5ecb906d5ea831724ed430013;
mem[90] = 144'h08c5ff9c0ecf0069fd37000f04faf872e5f8;
mem[91] = 144'hf8e3f4f10d900b8816131402e09bfd111dfa;
mem[92] = 144'hf01fe29eed59ec4af103181e0d1b0067e634;
mem[93] = 144'h1f4becd1095010ee0143f9dafe82f3440a63;
mem[94] = 144'hed7317a81c7f1255e47be71616501b171db4;
mem[95] = 144'h1fadf199fb28e137f0f5ed81e2c419171611;
mem[96] = 144'hec31e7a1efd7f180f9b50e8ff42d0a21fd06;
mem[97] = 144'h05a01ec71e7e0f1be077ecb40f57f160fac4;
mem[98] = 144'he842e4b705b407801ef8ee871026e894e5f6;
mem[99] = 144'hecd71f40e612144ae73314a70d120a0505ae;
mem[100] = 144'hff4eebed0b3ceba21e8ffa940076199e080e;
mem[101] = 144'h0233ee83e521104f13e30f780b5a0fbc1ff3;
mem[102] = 144'hf8cbf0541a581abce8cbe1a3f6910d600c9b;
mem[103] = 144'hfff417db094306a51949e17ce6f30df2fe30;
mem[104] = 144'h063c176cf179f4bde831f0721b9c1b2e14ab;
mem[105] = 144'h08d6097718c200c41514f62219deebc6fab2;
mem[106] = 144'he3110ddaeeabf63f135117f206b1f9fee5f6;
mem[107] = 144'h074b1fd20b86f9e20f56085a19141206e5e3;
mem[108] = 144'hfe761a970ae3fbb6f536f4501cc0e612eaa0;
mem[109] = 144'hfc22f24e05a0ff0809381b361470e2b6050f;
mem[110] = 144'hf99e0455fab7ff531140068ff241f97b0f4f;
mem[111] = 144'h0ff01b21ffc009f6038600d710c7f2671b84;
mem[112] = 144'h129c0a521677eec81ff909d619e500af15dc;
mem[113] = 144'h002f1db515341a0ee928f050193ce486fd3d;
mem[114] = 144'h1c8a1140feb3f6c11dbb0dae1946e89d0833;
mem[115] = 144'h07bde13a1a2c086518a0f5fa09b3f1c20fb6;
mem[116] = 144'hf22fe34df9981b56f021f4aa073500741818;
mem[117] = 144'h090bf0ace9550d3806c3f1d7f839e3e6f201;
mem[118] = 144'he2d80b071e17f58dfd4d0ba00d68f5480e5d;
mem[119] = 144'hed9feab4f8e91380190519f41837f2111ec5;
mem[120] = 144'hf5f61aebe385e640e208f927ee1eed8a051e;
mem[121] = 144'hf68412910c6408ec0c06fe69e4d50eafff3d;
mem[122] = 144'hf2b3fbee0c081ee6f82ff240125afe970649;
mem[123] = 144'h175c1e3a0950e80503c2e6270b1d1301f3d9;
mem[124] = 144'hf50cf6091a96fa18edf70c91f9d60421fc02;
mem[125] = 144'hed69ec76fa17e3bf1cfb11fefd07f6711558;
mem[126] = 144'he014edb2f51317d5fdc7ec0b0ae3fb71ef25;
mem[127] = 144'h17b21081e110eef505b9fd770b71018816fe;
mem[128] = 144'hf1af03fcff3001d717f71e7f14a81a710469;
mem[129] = 144'hf81cf442fbd40a58e45c12f1f6d306f91ec6;
mem[130] = 144'h18bb1455ecbdf73e0aa60e5e15e11395ec4c;
mem[131] = 144'h119af67ded57f77201fee8bff53e0d630909;
mem[132] = 144'hf1061c6b1be00db2f23716290bf115b0eb68;
mem[133] = 144'hf58bf88eea70fc5016e40dcffbceec301143;
mem[134] = 144'h1f2917060cd6ed6eee9e0f3a05af0775fc73;
mem[135] = 144'h136017521c59016ff2181264f5050464e5b9;
mem[136] = 144'hec431269e17800f5ee661e85e5cd154a1f50;
mem[137] = 144'h1eecedb8ef5de8afe2fbf66f177e109f1b18;
mem[138] = 144'h03241a3810d70b7903dcf17d173eedd611a5;
mem[139] = 144'h038e10781893fdf2f0a612f6185ff1e3ebaf;
mem[140] = 144'hf3a20855f7ddf340eea71b2018010529029c;
mem[141] = 144'h1ab702b7f0e6ead0149309faef0fec08e52f;
mem[142] = 144'h059c15af1066f0161d7415951607e79109b1;
mem[143] = 144'h12b8138af2371eaf1d20e0ec19c4e5c50695;
mem[144] = 144'h17befb831dc6f7e80954f01815fdf577ef80;
mem[145] = 144'h1e801eaf1277e8801068fa46f03f17091762;
mem[146] = 144'h00f60f63ef4ce4620e79f608e860019611ba;
mem[147] = 144'hefcc0238f87418cde05a0a9e0161e857003c;
mem[148] = 144'h10f5faebfe7b154615a61cabe55f04540951;
mem[149] = 144'h1edf180a02781495ea0be647021c0fc6e23f;
mem[150] = 144'h0179fe3eefbe04c70369e991e6f6fd5ff508;
mem[151] = 144'h04730a4a072ae678f404008c1ed2e67e06a3;
mem[152] = 144'he053f614070ae2e0e8bdf54602fcf893f00a;
mem[153] = 144'he8561db617fff0df0bc904ee1b071e8201fc;
mem[154] = 144'h19d7fd00f667ec1ff9cafe800264146116c1;
mem[155] = 144'hefc4e9ffe3221ce5e923115503c5174a0558;
mem[156] = 144'hebe21da4e2f2e60df82318eee44f00da139a;
mem[157] = 144'he6f7fdfee8d31fa5f198194bfe55f1c5eada;
mem[158] = 144'hea5b1b1d0352ee10fe27fba205621b11ea58;
mem[159] = 144'h0ee0f5550c301842170a08d5101416890358;
mem[160] = 144'he815fdd5f92ae62e0526fd31fba6051fe473;
mem[161] = 144'he8e6f05af9a50fb80a7a17fe07a4f2e01503;
mem[162] = 144'h0b7b108711ef1780f561e219ec1b1c6f1754;
mem[163] = 144'hf7a50fdc0a42f00fea6c1526e19601891c09;
mem[164] = 144'h05660627f9beffc613560eac0db411891895;
mem[165] = 144'h18b51d62fe03143af4b21a7ee353e6fd17a9;
mem[166] = 144'h15ff1a660b2f0298e487f3d50965ee0302cf;
mem[167] = 144'hf51ce6fe16340b6b0108104c05e61c8ae274;
mem[168] = 144'he885e46f1bdb00f010b103abfbb8115f0ff4;
mem[169] = 144'hf18cebce0e8e0dfa197a03e5196a0bb31249;
mem[170] = 144'h0d34fb70efb7efb40f6be639066e1bd014aa;
mem[171] = 144'h086213fee1d51905e352f9a7102c1ff4050d;
mem[172] = 144'hff14e0f8fdb9eee311db06591372fb0bf068;
mem[173] = 144'hff5ef6330da8129be94c091116fae912ec4f;
mem[174] = 144'h00d9f26df20201e5e3150edde44a0764e1a4;
mem[175] = 144'hf416e4ba1b520770fc53e9a3ef3d10c500a1;
mem[176] = 144'hf2841767ee39fc77e7fbe498f0fef6a9196a;
mem[177] = 144'h000cfc9012111368e574e5c219591ef5097d;
mem[178] = 144'h1e841d840782fd51017515fee9d51f41f559;
mem[179] = 144'hf5d51e151083e436f0c80b1ce16de2f006b8;
mem[180] = 144'h027800deec2a1da5f7ad0bc4f319f404f009;
mem[181] = 144'he6d4085df0fb143c0083123aeecf1e800f7f;
mem[182] = 144'h1914e3e7e594f82ae686f5450ec8fb71166a;
mem[183] = 144'h010b1e54eb6414631b42071bf09df75af2ba;
mem[184] = 144'h025910d80e0de26ee304114601d9edbff3ab;
mem[185] = 144'h0eb60c100e6e000ee3d71d8f0af51496e5f4;
mem[186] = 144'h1f1bffd1ee3ce63412a50bafe89a17b9f2d4;
mem[187] = 144'h00251e9be12ef1bef2c5ea0cec941355f11d;
mem[188] = 144'hffd9fa6a0d240ed30145e77df594fdbb0159;
mem[189] = 144'he371ed1bfcfdff9d1559fa200884f090ff97;
mem[190] = 144'h0226ffc4054ce4c9e785ec3b005df4b31766;
mem[191] = 144'h0a46f498fc9ee5241133e39e186315f3e12d;
mem[192] = 144'h0da21d2509531a901b4c1ae1115a0d46e7eb;
mem[193] = 144'h0aca1c0318e71331f5d9e649fca4f9581a5a;
mem[194] = 144'he808fddae939e4f8f17f114de1dafa3ce8ab;
mem[195] = 144'hfd350c7deb130e89e27de8ed131be67c08e4;
mem[196] = 144'h1f671955f59215f9f738090deeede6e30585;
mem[197] = 144'h07b3f1d50b2c0011f92be9b7fb45117ee6fe;
mem[198] = 144'h0be1ff341df3e57ef4c1ebf1174208e51a76;
mem[199] = 144'hfa75ed141a69f8110230fb05f68c08a5ff0f;
mem[200] = 144'hea0d0614e30ef860ed7403401950188be153;
mem[201] = 144'hfd58182f0a0fea55e63dfefef853ea50e671;
mem[202] = 144'hf92afe45efcb093509c31883e950fe980be2;
mem[203] = 144'he89bf9a6faf1f35df956ef571d35e986e862;
mem[204] = 144'hf2df18f81b970e42e8e9e8dc11a1ea91ee9f;
mem[205] = 144'hf6e0f815161c0f5c0484f1d31955f73ff376;
mem[206] = 144'h1169fb71188cfaa8edb6ecb500be0392ea52;
mem[207] = 144'he117e030104812520326e055ea8bfeb8ef1b;
mem[208] = 144'h10c5e566fccef67ef3f31fc7083b0e0f02be;
mem[209] = 144'h1695f544f4fd1196f5b6f06308661657e072;
mem[210] = 144'h1025125e0dd319e80df9009ee095f7c110fb;
mem[211] = 144'heaeff17d011611090b9df83be6e6fe020cf4;
mem[212] = 144'h113aebe4fc39e74af164f437f4510c72ff29;
mem[213] = 144'h17c1e5f4e7f8ea78f1f3faeee9231fa2176e;
mem[214] = 144'h01241a8c0a8efac4081e0bf5e172151b07ef;
mem[215] = 144'h02c002bdea67e0010b7eefc8ff321dd3ead1;
mem[216] = 144'hfb5e041a1722055d1e61f26ce479fc90f192;
mem[217] = 144'h16361d790d20f733f974fe5cedffe4a4f148;
mem[218] = 144'h0402098d0ebf1e3c1f0d1aecfe191e65e801;
mem[219] = 144'hedc7e7111234ec74048af7efe15f038a0ae8;
mem[220] = 144'h13ca17f1edf1e6e70870f65be3f4fe4a151f;
mem[221] = 144'hee79e393e272e92ffac0e0990f500119f840;
mem[222] = 144'hf92e01a9f587141d12a5efd5e978eec7124c;
mem[223] = 144'hf6e518d5050b1c98edbbe0c315280ff7e5de;
mem[224] = 144'h0d5d01ddeb8e04fd1bc5f953ed780fe5e28a;
mem[225] = 144'h1c820143e09eeb6f000ce2bf00baf4dff1cf;
mem[226] = 144'h14eefb0bf9b2f20711cb0d3f062cee85f464;
mem[227] = 144'h0fb81cdf1fb4197ee1ce0b6a0c150d7b171a;
mem[228] = 144'h0583e5fce8d51beaf09b0edbf20d0f7915b4;
mem[229] = 144'h05afecf2f01d056118dd1d1c1f3df44e1494;
mem[230] = 144'hfc49ff59e73e090b101c0423e9ad0d5c011a;
mem[231] = 144'h1e0ce139e867e10be733ed34f1b5023206f9;
mem[232] = 144'h1afb0bc9e3381be4f135fee4e4f0193b1f74;
mem[233] = 144'h1f2ffcade049e7ba193c03c5f7f7fe941ca3;
mem[234] = 144'hf28bfe51137b0b331ee61da80e71ebdc09c0;
mem[235] = 144'hec35033f1cd6f9291f03f5e8e581f283eede;
mem[236] = 144'h0e6113deef8bf9cd10fde4ab04d3f98e172e;
mem[237] = 144'h1234e012f334e2a017d3ed83f7e7f8b3079d;
mem[238] = 144'he6f91e98f1b51bafef10e0c60fc7ea4ae56e;
mem[239] = 144'h0421f704e7cee4b906c5f148e0a2f3641354;
mem[240] = 144'h0c66e4c9ea21e806fc3be191fd8606b00514;
mem[241] = 144'h15850722e99afc5de532e4acf1ff1df4e032;
mem[242] = 144'h12031c66fd98074ae53012a306fbfc8cf027;
mem[243] = 144'he6451a170d4a1114ffff0105119a067cf84c;
mem[244] = 144'h129de39f1ebe0c0e1fa4ea17f009f967e34f;
mem[245] = 144'h10ff0f9705b51a2ff394ec2116470ef9e03e;
mem[246] = 144'hf854feffe54ce80efc8c02d4019deb82025e;
mem[247] = 144'he4ca050af1b1f09c06d2f4b41355e217004c;
mem[248] = 144'h14ed08111408e116f8b40a97ec9ef6fef83e;
mem[249] = 144'h17eb0a4015730e090aeb0cc3055cf75b1e6f;
mem[250] = 144'hef5b000311b802fffca7174a0f9306d2f176;
mem[251] = 144'h03ce08cdfc8d1dd3f18cefcf0408182de28e;
mem[252] = 144'heaeefd8ef12c1e58fcfdffa803401fff04d4;
mem[253] = 144'hf8e4ed55e525e9a9e0f7fd2b0943fb74e90d;
mem[254] = 144'h0cc21961e4681d031b06fc761b39e4a2ef4d;
mem[255] = 144'h0c7de9841050e7abe7b80e01e1e7f100eeb2;
mem[256] = 144'h1995142a07a6e7f90baa17d90fbee96509d9;
mem[257] = 144'h0109f5b20e10140702b5f61103620741e8e8;
mem[258] = 144'hec37e0160d440a5cee2ef52a1ad0f10aecce;
mem[259] = 144'h18fafd46e5281c9afec41e9812a8ed1d0d93;
mem[260] = 144'h0322e30cfc23f3a8e2f610a5e7e8f62e0f54;
mem[261] = 144'h0fdc0ba1f678f28914eff1801b6614310a41;
mem[262] = 144'he20af18ae2450bb6eec81bbfee80050aea22;
mem[263] = 144'he305fbe4f62b1c56f1e6f6d6f105f5601248;
mem[264] = 144'h1f1d0f72f3b5f404e3e01ce208fd0c701f79;
mem[265] = 144'hf9ddeb6307caf17214c4199befac09c40e2c;
mem[266] = 144'h0dcb0783ea6405dc1ebe196ef631fd481d3b;
mem[267] = 144'h108212a1e64c04ec1fe5f144e1cd10cce298;
mem[268] = 144'hf3c7eef7eb94194f0925e4331328edd61d88;
mem[269] = 144'heae20b33ecea104114d712e3e483f749f1cd;
mem[270] = 144'hfe841d6e0b9401f0f9440354e9c11c3eeb52;
mem[271] = 144'hfe7ff97bf8dd0cc307491148f7c4efce1140;
mem[272] = 144'h0d3ae0b8fbc1fee80ee7f43e106ff653eb56;
mem[273] = 144'h1d2a05ddff0df74bf4df0eb905701aee02a5;
mem[274] = 144'hfb6f1ecdf9adeccced0d1a7a0ef3fd62e46a;
mem[275] = 144'he5410eece2c20242f1cdf1210d68079a0180;
mem[276] = 144'he4e40bb1137217150b49e5e20ac3e37a037d;
mem[277] = 144'he81501e20175f69deb86e36f17d6fa960861;
mem[278] = 144'hedd1e5c9046414c003d4e1fe15dd11b1e888;
mem[279] = 144'hf199ec46e5a9f9a8e762fa1cec2be551e8d7;
mem[280] = 144'h16cb0e71180e0a1eed231a18f47f058ef099;
mem[281] = 144'hf3c8047ef2d80b501761f2031bda12000a99;
mem[282] = 144'h01180f0ef6300cf21621ff54e3baec84fa91;
mem[283] = 144'h0a63e3bc1c60e0bc060fee7a059910251d47;
mem[284] = 144'h0c0a0979f9651fbf174f0e6ef838f49df969;
mem[285] = 144'h0ecdfba1e753f136ed2ae6cd1418fa4af227;
mem[286] = 144'h1c38ee7de69adfe4013afaeff6cf082416b3;
mem[287] = 144'h10eee9751d53ea22e27fe0ff0845e8a6099f;
mem[288] = 144'h1239f13d08ce120d16ef16dd0380e190fffb;
mem[289] = 144'h08a4ee48022b1380e70203e41b62f76beb52;
mem[290] = 144'he0ed047ee0ec1d7007f104e9f346fbb50353;
mem[291] = 144'h120403baff6f1d6c05ca177b1c940cbff744;
mem[292] = 144'hfe5bfe6f14551cb4001c1deef1d1f7fefb7d;
mem[293] = 144'h08c01599f574f51b1678e980f941fc96ed77;
mem[294] = 144'he5760a9e15aa169eed970a63fb86108f05fe;
mem[295] = 144'h077f1b8dec4be99917e300ec0f91126ff608;
mem[296] = 144'hecdff5880165f5321601164ce698145d0993;
mem[297] = 144'h05b2180603b50b5108580cfdfad707e71750;
mem[298] = 144'he1a3fe62e1f7e76be247eec9faabf382054b;
mem[299] = 144'h0d7df79218b71ae7feeee1b917d31cc0f942;
mem[300] = 144'hf69cebebe616f97deac00f8f0231f2041843;
mem[301] = 144'he24f1edfed18ea0ce9630b55e3ec13b2fb5a;
mem[302] = 144'he9c7e7ec15c5f62ff8d20ab3f24af7f5f8b7;
mem[303] = 144'h0e7ce3f3e3781d930e62fd9bffaafb98f7bc;
mem[304] = 144'hf5420d980537ff3dee56167c1500f4bae061;
mem[305] = 144'hf065f65217df13dae8240a7af693e114e42f;
mem[306] = 144'hf4d2f62de4c70a970e6af26dffb8f09ef9d8;
mem[307] = 144'h16511f9cfc971e9bf262f7ecf313f426fbd2;
mem[308] = 144'h16621b54eed20ba3e74006f9efd8f77b11e7;
mem[309] = 144'h19d4fdd8e1820ea8f30be525f82104e0fbba;
mem[310] = 144'h1300e8041129067ff16e119cf32aefde069a;
mem[311] = 144'hf97013b3f4e1f3850ad41a2b0b85f9dae960;
mem[312] = 144'hf4def073feaef5cd078e110603dfea880dfb;
mem[313] = 144'h134fec18e720f0d904e507db09a5e2bffb9a;
mem[314] = 144'h19f812a2e235e628fb0ef7f6fe53f4570ce9;
mem[315] = 144'h02e4189cfd8ef0631e59e5dc199904800411;
mem[316] = 144'he8b8eda2e93ce6f4079afb1a1ccbf129e267;
mem[317] = 144'h012b1faf1c38f181fa68eab51431e97d1a7a;
mem[318] = 144'he13a0ae404a5eb6d0e02f2110386117804e2;
mem[319] = 144'hf6f9e01c17e80aa9f55e1220e50d19b919dd;
mem[320] = 144'hec3218b7e259089b1b2e0c1cec37024f0aeb;
mem[321] = 144'h12491359e50f1747f9d5ebc2f62a00cf12ec;
mem[322] = 144'he89f03ae05d302a41566f114f086e88e1000;
mem[323] = 144'hfcdbf8eaff2301641adbe8bd1fbb13810bfd;
mem[324] = 144'hf9ccfa53090a040bfd8619470466f22ff963;
mem[325] = 144'hf55cf4a2f9b50cace1f80d87e1a610cf1bb1;
mem[326] = 144'hf9b7e6f11fe81348eb31097304f0f5f3092e;
mem[327] = 144'h0d3d0ab7115fea9be93ae77c0cdbe857ff42;
mem[328] = 144'h15f4eee4fce412440ee8e87ffb6eea9f0dd8;
mem[329] = 144'h06f40152ee3bfedcfd45f256e2ea0371f09f;
mem[330] = 144'hee140168feb307f81d4eebd2e3a306baf268;
mem[331] = 144'h03db0c3aff1dfce51ceae5840665e68be007;
mem[332] = 144'hea51e8c918431c34049cfc9ae7c00aa4f367;
mem[333] = 144'hf7bee4d1f132e6b615d5fe1b1d560cd60585;
mem[334] = 144'h134e15390ba0fffb1b1a18ecfa0fe4410b7b;
mem[335] = 144'hf3e106091529fb8e115df58e1129f95e141d;
mem[336] = 144'hfe640f921080f3391e7119ebfe15e3ae0402;
mem[337] = 144'he600f913e073ebfdf5cbf69ae76e190b096a;
mem[338] = 144'hfcd5f330fc8b179de13618f90ee7fad5ff2e;
mem[339] = 144'h06be186dea9e161ae063e54b037ceb65ee85;
mem[340] = 144'hef2817aef080e9990dfeec6de3491a85f6dd;
mem[341] = 144'hff6b0596004df1d7f7bee47b1195079dfd44;
mem[342] = 144'he330fc5806b80e6611a31f06f6100ec4e40d;
mem[343] = 144'hf8ccf3431a13f7f211efeb86ea7f0d5afe12;
mem[344] = 144'he4501badf5bbee97e8fe0a510d71041e0f1e;
mem[345] = 144'h1760fa6d0247fee1fc501a26f64114c5fb50;
mem[346] = 144'hf12a1f80e18a18b013c7f5570831fdc8e896;
mem[347] = 144'hf4d6046b0a7ff5d8fc3c1c161a180625e0b7;
mem[348] = 144'h0ce71fcef636f852ea45063cf71ff085f76d;
mem[349] = 144'h101effa5e9d7e6bc1473e378057b117507a3;
mem[350] = 144'he6aded5800500a220ac8143d1ac81c02f571;
mem[351] = 144'h0c8ae7b016510cbb1c641158fd4c1755005f;
mem[352] = 144'h1378ffac04a31e9eeccb17e21e55fca71e53;
mem[353] = 144'h0b27091108e60425f31ce8ef10e4e6111b3a;
mem[354] = 144'h04a0ea2e1b4e03a7eceff76ee7790070f8a0;
mem[355] = 144'hf6b0192bf715197904210f4909fdef721ea8;
mem[356] = 144'h02a80d71e7f11f1e1d7b1f3c14af0a400a35;
mem[357] = 144'hee6d08eee84b1783f8b1018cf68af425e6fe;
mem[358] = 144'hf4410365f77a0ceae5431d1f16d9f262e3eb;
mem[359] = 144'he812e3adf6850a86f8e8fe0af8b10a6015db;
mem[360] = 144'h1303fc90f943e4051f1906220a1504a6e70e;
mem[361] = 144'h1ca5f909065ffa0be59b1243f2d90193169d;
mem[362] = 144'h138c09d1181ee8c5f32b0172f837f7be1726;
mem[363] = 144'h1dd91c201a5ef918f54a06670f481bd9ee61;
mem[364] = 144'h1da4144a1837ec6f1258f2b0e93a064fe668;
mem[365] = 144'hf16b1ed009f801511f8f08d3ecbb1b94063e;
mem[366] = 144'hffe10b1ce3f2e0a3ff090f67fa5c198c1af6;
mem[367] = 144'hfa44e172f2961ca91086fac7ed591566f0e1;
mem[368] = 144'hf410ec80e3a71e3febaa15c501a6e9bee6e7;
mem[369] = 144'h0649f92415deff97179411f609ee0180f080;
mem[370] = 144'h12b10a94e613e15ffe06e99a0fbff4c2e3ee;
mem[371] = 144'h1095f8b4185e1b99f799f7d01c8106101e71;
mem[372] = 144'hf79c1c50fa0d142901d9ef72e25dfb3cf93a;
mem[373] = 144'h10e6e11e073be57616d111cdecad134d0b79;
mem[374] = 144'h17c21d9be11c1c160311100af257fc7b06c4;
mem[375] = 144'hf6c9e47ef8da0ed4f427f3fa08abf1d70219;
mem[376] = 144'h0d85108df8f01bf10afefb9d1cca17fae8b0;
mem[377] = 144'hf4b9fd7f18bc17a0e1de1bf0f3b91e641339;
mem[378] = 144'he41502450b6a09e8ee77127ff5271c13f3ad;
mem[379] = 144'he742f398007bf32dffcc0aa20c141db01f15;
mem[380] = 144'h165509eef524fd2ef8e80a7e05ae0ca5e923;
mem[381] = 144'he6950486fa98ed400b13ef4c03691afee10d;
mem[382] = 144'he25515d216590871127a10a4f54ffe700f2e;
mem[383] = 144'h1cae056618feee8cfe6617ddfd8604b600a0;
mem[384] = 144'hf48bf418ee76ea3c176b1352f5320dfde39e;
mem[385] = 144'heb70e93e0ade07d71ce301eeed140594e801;
mem[386] = 144'hfadd0bcaf807fee5f8381c9113d40bd2edae;
mem[387] = 144'h05b90e910fa8fd4df7c5f85bee611793f28f;
mem[388] = 144'h108cfebbe4551a621bdeee4df1190802eb6c;
mem[389] = 144'hf9e8e25a1da9e47d1b14e4910c1f10d91e0f;
mem[390] = 144'h1b9c0490ef0eebf90e99e624fc3c15d6fa18;
mem[391] = 144'h15a40b02ea29e8a417201bb7e9cbff991459;
mem[392] = 144'hf6d8fa5905f6e3ca19270e61038c06480597;
mem[393] = 144'h1de215e2e9a5182713e41914e6d0021c1917;
mem[394] = 144'hec7d1199146d13faeb62069b07fd1a6b15d5;
mem[395] = 144'h0adf132a0feae20e04e0111e105d09faf70c;
mem[396] = 144'hf6c405b31446e75616b7e70502f3fb8ee902;
mem[397] = 144'hf80bf68706cee76ce606ed9ff5960a3deedb;
mem[398] = 144'hffdc1d9d01edf281e04cfc200da3e5a3f74b;
mem[399] = 144'he4c6fcbc02e7e3390ac013381ce604a4f598;
mem[400] = 144'he95af55de065e66611c503a0f06d0d0607f8;
mem[401] = 144'h023ef8d9ecfa13d6fe7afa4d00a0f984e72e;
mem[402] = 144'h021512b702f113b5f5c909a70fb2fc5b02cc;
mem[403] = 144'h07241a68faa8108de153f3551ed11462f5a4;
mem[404] = 144'h1138fbd0e7060bc61f55f9baf3570668e37a;
mem[405] = 144'h1d72e387e5bd1df7f0670a4fed92efbafbd7;
mem[406] = 144'hfb3fe4d70b7719d509d2fe2411041eb9fbf6;
mem[407] = 144'h0e0402e41634efe61a92182dea730f7d105c;
mem[408] = 144'hfa390d52e5f1e3ccefa11d78e609000f00e6;
mem[409] = 144'h0148e6c11fb3f7560b27f57c16f01c40e8b9;
mem[410] = 144'hfb87f9d1ec810325f8c1e432f53f1dd702b6;
mem[411] = 144'h1870f918ec5602801da40b1a12851685e5e0;
mem[412] = 144'h06a805f31af0f60a186ee6ecf578e2081b1b;
mem[413] = 144'h0d0ef6afe8fc112fea5901fee9ca0be1e0e2;
mem[414] = 144'h16ad11a5f239e2e41a070602f52c0e5dea9a;
mem[415] = 144'hec441ace1847e22b0f8e08091979f6c5e625;
mem[416] = 144'h0a91eb47070af32904d610281dc00969e199;
mem[417] = 144'h0fc81ed20a7a0fcd02e1ebcc036d05f6e299;
mem[418] = 144'h1b3ff650e7260f1be4161eddf594fbe2fa48;
mem[419] = 144'h15f719dd1a121c150bfcf2daeaeb05c41fc6;
mem[420] = 144'hf62a00c601e4f365fdce11fa0a631ec1efd1;
mem[421] = 144'h0731e418f3c108010503fbd5e723007aef3b;
mem[422] = 144'h176ff733fb751b1a09cbe6aaf8830755e515;
mem[423] = 144'h0444ff0aeda31e7df16e1f5213ecfe07e27f;
mem[424] = 144'he43a0ab3f92201680771e3f3fb79f37108a6;
mem[425] = 144'h0ee9055dee64056df1d7079fe1b1115b118c;
mem[426] = 144'he1aae1cafd40fa7aefb60b5b199904cfea34;
mem[427] = 144'h0f371c7c0f271a9d1dea04ff13fd01d30a0a;
mem[428] = 144'h173ffb95e2cc17f9035def71f2da00ef1075;
mem[429] = 144'h05f5fbca131318b518d8e39ceb5fed52e5b9;
mem[430] = 144'he572e7e70da0f049e943e41b02a9e3f80184;
mem[431] = 144'h07a2f5d6f7f0f94bf64007adfb03183be0dd;
mem[432] = 144'h08741f8f0cdb0db516941a970cf2e2570278;
mem[433] = 144'hedd81b7df1bdfadbec811ad2e67cf2940a02;
mem[434] = 144'h198bf00119e204a110baec68056612c119a9;
mem[435] = 144'hfd3fe536e60813de037df0a11c3ae025127e;
mem[436] = 144'h1deb0191ed890ed6f74815b6080c10eb19b7;
mem[437] = 144'hf6a1e49101df114af4f1f93a1c51e96918cb;
mem[438] = 144'hfec3e13fea840e3e0c0bf7d1ef48eb4cf9e5;
mem[439] = 144'hf1e6041de0080d0c16afec7114aa18c9e6ac;
mem[440] = 144'h158f1a9419511e75fb31f188f3d7f72f1a55;
mem[441] = 144'h0960fabb1d38138cec55fdcbe85f1f42f393;
mem[442] = 144'h090816fdfcb5f1c5ffdee3611289fb6ef956;
mem[443] = 144'h1c0af0810252f2351eefff9109eae9051444;
mem[444] = 144'h148301c40e3ded230cb9f7ac047eec62157f;
mem[445] = 144'h19dcf964119be874e543fdea1b64fa7c0c3c;
mem[446] = 144'hf6e20527e56f00f11080f339ee84e7e1ed4f;
mem[447] = 144'hed8be1570ed0028d194ffeefeae1f511e3d7;
mem[448] = 144'hf71108bafb511a4710a9f9e50a2917bc01d3;
mem[449] = 144'h05ed0c75ed15fa7503340c291ec8fe83f02a;
mem[450] = 144'h02dff6150888e093f9c5150afe031432e39a;
mem[451] = 144'h1880e222eb9b1b8b10fdfda91d3f1c7312e0;
mem[452] = 144'hf6c6fe05e1a9f1ade5c8fa350d970e021ee0;
mem[453] = 144'hed571dbffca2e94efe5f06ae16bbe84d1cfa;
mem[454] = 144'h1a22fdb102bcf7c9e70fe477f936e41ae732;
mem[455] = 144'h057613c31d8afb5ee43d1471182af6fff28f;
mem[456] = 144'hf3020f380009e309f8b7044c0eb314eff6ec;
mem[457] = 144'h0be6f24ceaad0fd2f934e7c4133f02b3ecd6;
mem[458] = 144'he1a117d1eea60b1efa11f06fe194e05ae49b;
mem[459] = 144'hfdd50464e89a1a5dfc12f170037210a5e999;
mem[460] = 144'h16d5f51f1f1de2771fefe6a9135a08220d16;
mem[461] = 144'he5921017ea980febe691e29610c3e6ae03bb;
mem[462] = 144'hfb2cf571f012fd8ee047f6090c1ee9fcfc76;
mem[463] = 144'h0435f2de0298f22ce1cff952eb47f93212a7;
mem[464] = 144'hfa720c811ebc1deee63be5c5fb44fd48fdbc;
mem[465] = 144'h08a601f3015d04f3ea77140c0d7ee7230391;
mem[466] = 144'h19acf50919f30df90b28ff9ae5961023fc63;
mem[467] = 144'hff9704a31c97fc9912a51f3aeb3412b8087a;
mem[468] = 144'hec5d1d591fa007601607f9c1f1a7185dfefc;
mem[469] = 144'he4e9e5521c29f4170f901fc417380a49f8fa;
mem[470] = 144'hf0091d27058d0cacf6a91a52ec890bd91f7d;
mem[471] = 144'hf8e712e91e79e9340898074fe79d109502dc;
mem[472] = 144'h1967f4661a72fcf8198a117feca00164fb61;
mem[473] = 144'hf7bb16960a85ed02087c1be7faaa0c77fad3;
mem[474] = 144'h047c1b8de71306cd12d71f4e163de19ee916;
mem[475] = 144'hf1d517ee01f50681152309a000c90ccd190f;
mem[476] = 144'hfeacef6bf50ef91cf25feb44f97df3cf0dba;
mem[477] = 144'hfd89f1d6efa4fcf3fd6d1848106512440401;
mem[478] = 144'he0761765ea031405ea45e90ee690fca80a26;
mem[479] = 144'h1dbaf726104017b40b49ffdd02ff076ae056;
mem[480] = 144'hf6aee6e413fefdfce53f1be9185611fc0163;
mem[481] = 144'hfab70c16e832fda71d7af96de87be7e5f055;
mem[482] = 144'he3511b5c0859fcbf034305cf150a1283026b;
mem[483] = 144'h07dde098e6711557efbff8a3e37af98e13f1;
mem[484] = 144'he5d416ca0fa8f2dffa7a11641fc0e0aee943;
mem[485] = 144'h0575fd230e26e0090acfe828e80ee4af10d9;
mem[486] = 144'h01b41e9213ebeb62060e064ffc36ef130d91;
mem[487] = 144'heb16e72e12befd59183def0e0908e49de776;
mem[488] = 144'hf39d18d2ea3412a81607eea0ea0e041212cd;
mem[489] = 144'h0d60f4a8f564ebbfee2a01ce1d34fe30e336;
mem[490] = 144'hf4f2068f05780837040f13b304f706370805;
mem[491] = 144'hfe9f0b9506f9e84f00bff87501dcf20200a0;
mem[492] = 144'h0c5e1675fab4e0c20d70f01e0c16eeca1cc7;
mem[493] = 144'hf7f815ca140f0e81f0991cbfffbaff16e042;
mem[494] = 144'h08ae15cd1a2ff95be1b40d68f72ce6c81e2f;
mem[495] = 144'hf9b41257e359f9f4e8fa1ec317e81279ecd6;
mem[496] = 144'he669024cf6d2f146fb95056b080e113505bf;
mem[497] = 144'h0c05e469fb9605c6ea4dea38ec8a11c00593;
mem[498] = 144'h13c01064e0e90a37e34be2df0be70015e894;
mem[499] = 144'h03fbecb1f8d51f37ecc91c5ef12a17e7fcae;
mem[500] = 144'hf40cf38e1edd012b1079eff2f33b049400bf;
mem[501] = 144'hf0e11d320f3903cee417ecaceeb0ece7e667;
mem[502] = 144'hefabe927fe381c24f6411ecb07940a8afdd1;
mem[503] = 144'he18d0011ebd4066be77912b203ffe0b106c3;
mem[504] = 144'hfa05f291f2c4156a02e5ffc8ee8a0fc2f2fa;
mem[505] = 144'h0337e30800d9efc3e28d1a6001c7f04ef230;
mem[506] = 144'h1eedecdd050be98408b7eff4e5f4e871e322;
mem[507] = 144'h18aeeff6fd14e1100533ed90e011fcc70f3b;
mem[508] = 144'hebca1a8019eaf540f948190b1a28e5ac08e9;
mem[509] = 144'hffec11d1189c101aecd4e285ea13fbd808f8;
mem[510] = 144'hf56df3d7e004f2cdf4d3e723e22414cee0cb;
mem[511] = 144'h1240e74de3ab1511020fe44cec18f96be905;
mem[512] = 144'hf3cd0946e321e3ed1390eef4025004871fce;
mem[513] = 144'h05e81e1c116ef75b0038195bf3d909f60674;
mem[514] = 144'hf56ff272f43d1034f3ae0420f11c0388029e;
mem[515] = 144'h0e30e152f278f79ef774eaad02f20b281525;
mem[516] = 144'h1d550e191ce30f4a0375176800141e2f1f96;
mem[517] = 144'h055c008d08e71b0219ba18cc160a1670ee4f;
mem[518] = 144'h15a9f1591a82ee5614171a64eed215e1e715;
mem[519] = 144'h1a89e477e98a10451afbfbbc16d9057009fa;
mem[520] = 144'h16d51ac71582eba11322eda5ed640a0605d0;
mem[521] = 144'hfd000f27fd8017dfe5bcef3d1f4eeaebe5aa;
mem[522] = 144'h0c1df0b70f78e380e846fa180e5f1bf7e6ae;
mem[523] = 144'h0fad05acf3f80f49fd50e0c2f44715e5fe66;
mem[524] = 144'hea3ef82cfd6ef5a00cce0f37e741e45eeb37;
mem[525] = 144'h1d040442f9ed0fafefb0177c0857052e07bd;
mem[526] = 144'hf20d14640ce80b2416411a251c3c17b5156f;
mem[527] = 144'hfba7f683f3751ecd0838e81ee1a7eb43ee58;
mem[528] = 144'he50cf091184c02f3ee61f6050e1503f41877;
mem[529] = 144'he399139dfc79024e064c08c712790720e311;
mem[530] = 144'heea306cbe72813801dca088c1e0c085e16df;
mem[531] = 144'h02fe12b4e4aceaec0e0c1b33119def83e81b;
mem[532] = 144'h08dc16b2fe2f0f9efe7b0ba9e878022710ce;
mem[533] = 144'he25ded76e242fc7f0e22e3d913a30621e68f;
mem[534] = 144'h01a51e2017380684e788000417c50f20102d;
mem[535] = 144'h1629177cf08cebeb06b6e84d0fda16d8f713;
mem[536] = 144'hfe821f2c1252fa5ae6221e3ff96b1f641556;
mem[537] = 144'h0d1ae1ab0a4efbb2f4b0f4ae1d3018e0e2b6;
mem[538] = 144'hee71e6c01173e81afb0feb72fd38f3dfecea;
mem[539] = 144'hf5bef7fbffd4e2c9fe441dc2f83df689fdbe;
mem[540] = 144'h1fadf86ae2e1e4390e91fecce752f16e16b3;
mem[541] = 144'h003d1825054a11520bb5083d116a0606052e;
mem[542] = 144'hf33203d4f879e496123017fafc2f0be70b8e;
mem[543] = 144'h0f53eb37fef4e74fe2e31090f8891f06f5b8;
mem[544] = 144'he1d2148906f80423091a009214c8e089ea2f;
mem[545] = 144'h0e4a12fbfd38e4ca149ef00d0104f1521810;
mem[546] = 144'h14a211070849e1de1b9dffe1ebc3e645ecac;
mem[547] = 144'h1234ec37ec7514afe806104706a4eac800d9;
mem[548] = 144'hed52f3b11f34f9d2f1101e8e1972e4041dd3;
mem[549] = 144'h19601fe70910f65afc5fe554f1b20b59e15e;
mem[550] = 144'hf66311670165e1b3fa9ee3080ed019851da6;
mem[551] = 144'h17bb183e077014ace2e2047fe1f9051af10f;
mem[552] = 144'h0040fdb31b0b19a3f5fcf2ffe0360c09e596;
mem[553] = 144'h0e3ce062e81cf2f306d9091804c70d19f3a4;
mem[554] = 144'hf498e5f901c4f9b0fa640d66ffb21533038a;
mem[555] = 144'he40c1f7203e6eeaee73d076e187a1d8f1c69;
mem[556] = 144'he43b0192f1c71b69e15a067e083607f80c0d;
mem[557] = 144'h0cb5e794f4311013098d11be0db1e5fd1072;
mem[558] = 144'hedf00c2bfba5163afec21e3deb9d12a512d7;
mem[559] = 144'he7831489e3001b21e9d1144be23a118b1de1;
mem[560] = 144'hf0120135e442fe19f39f11d0f09f1f6cfaa9;
mem[561] = 144'h144b1c3a0392f6e6f8af0f5cef0dfe630650;
mem[562] = 144'hf6491627e3e311e9f832e3d1f332efb9e9f6;
mem[563] = 144'hfc911ceffab80593fb8416d3f43b171d0dd2;
mem[564] = 144'hf552ea091696ea4de8a8ebe0ef3b04241b83;
mem[565] = 144'heb381e13f46400d6eb08057ff3eb1dc20116;
mem[566] = 144'hf07506c701db11fc12e00c6df47aefa2177c;
mem[567] = 144'h102619091c71eea5e239e82e16a11d0218e4;
mem[568] = 144'h0ba31680ed8ff93602960be6093906150599;
mem[569] = 144'hec08fb3d02ccfbc8fb66f8f7f4aee5a21527;
mem[570] = 144'hf6fb0ddcf6eb017fef02176beb70e2230319;
mem[571] = 144'h08ce0d9e192beb23f8f611cf1da8eb0bea2a;
mem[572] = 144'h1f87edecfdc505d505bee0f2e7d8f120f243;
mem[573] = 144'h145616d90ec00ed7f8bcfe021b131f3fe88b;
mem[574] = 144'hfb4f0783e29cf4d3f8f30290177eeb34fe7d;
mem[575] = 144'hffe51754e736162401dcecf0f068025bf99c;
mem[576] = 144'hf6e8e11feeacf3ad03a0e995eb63f6830a03;
mem[577] = 144'he7361bb0178a0845106ae7d1e8aaef2104b8;
mem[578] = 144'hea9719ba0b230450078800f8fa510768e3ee;
mem[579] = 144'h1a5d114cf2c01d8be10c068efbbcf4e8efe2;
mem[580] = 144'hf5f4e4eff3c8e16fe4f9edd6e44bee9aef23;
mem[581] = 144'h0e240b15e678e5b7fa9fe26ef85c138df08f;
mem[582] = 144'heace15ea0b80f325181ee4be13f4188b1845;
mem[583] = 144'h072c08c5fd0919fbe81fedf3fe00f5a5f802;
mem[584] = 144'hf1d8f567f6cc059ffc74f7bd0383107612ad;
mem[585] = 144'h1901e751e87a059a1983e3611aa20a51e0b3;
mem[586] = 144'h150cee88f5c0ecb7f571f62c14651706fa7c;
mem[587] = 144'h1bf8e3c0eb49ff0efb7dfd14f05ff8ea0da0;
mem[588] = 144'hedee1d6df88a0de0fc2aede60c8f17370dba;
mem[589] = 144'hf38d1a8701a5f8f81ec01e1b08b5095afd46;
mem[590] = 144'he68a19fb0bf9e102fa7408dd053a03dc1294;
mem[591] = 144'hf4971a461b8be5c40c501ed90764f6aa03bf;
mem[592] = 144'h18d2eb6a093de9b118a502cb143d10db006d;
mem[593] = 144'hf66616360516001b0e430ff61865e688eada;
mem[594] = 144'he1cd0621fe91e4e40402e368ef23f3850a51;
mem[595] = 144'he58b14440cf6ff65e497e6e315f0f4d0020d;
mem[596] = 144'h19450fe11ceae6c7162ff407f767fc35e63e;
mem[597] = 144'he797e4e6e52f10ece037e6a5fac81013e230;
mem[598] = 144'h065a0b730bf8f74ff6e4020cfd5fe2d9eb14;
mem[599] = 144'hece10cdbf20c1d071762fdf2ff1ef45f0b5f;
mem[600] = 144'h1486e5590c58f4e6e652f8ba1ada04b8e3ea;
mem[601] = 144'hef43e716fac70db501be128d15571a3b169c;
mem[602] = 144'hf34012b019cdfe0506d5f2f212eb19f0f881;
mem[603] = 144'h1155fcacf8420e6bee5efbeb19ff13bd0335;
mem[604] = 144'h18aeec0ff4030e280564f7d6e68519c81353;
mem[605] = 144'h0c47eef00ca61fe9ed0e0f69fde0f734e461;
mem[606] = 144'h0211ed481387f8ec17ab1f90e362e9e409e0;
mem[607] = 144'he55c0e430892e0641ef70e221ec302b4e2ca;
mem[608] = 144'h0a81f5e4f78bfda3f892f8a01913ee9ce20b;
mem[609] = 144'he460e354f8d806381e720520ed5b1ca6e0cc;
mem[610] = 144'h1d25e463f38df01a152815feec7c1116e131;
mem[611] = 144'h1feffb44ef54f02b0d71fd250813f99cf876;
mem[612] = 144'h00440230e7461ba6f59210211f4ce654fa3a;
mem[613] = 144'hfe84ed8c19bdf8db02faf98ae43813190fed;
mem[614] = 144'h13e71b16ebb4e91213cf08580b43ff85f203;
mem[615] = 144'hf074f972e0c10019018bff5801030f40f492;
mem[616] = 144'h1fdd1fc91b97f1a1072ff855022d1306f312;
mem[617] = 144'hea26066d0846eb6515240abbf1430ef6f5be;
mem[618] = 144'h062cf43a0b121069fffcee24f4bcec1af37e;
mem[619] = 144'h19750ffa12f80371f7d9192cf7d3f3acefb9;
mem[620] = 144'hf59506a803bee3b6f2870ccdff74fe22f077;
mem[621] = 144'h00f91d18fd2ae1f509220950e9fc10140fbe;
mem[622] = 144'h0327e462004d0d74fbd3029118c50aff02b7;
mem[623] = 144'hfd28036603dff1ece392e000eb74e7790ece;
mem[624] = 144'h0c8be7c30347164c11aeea52e9bbfafb190b;
mem[625] = 144'hf37be5960a8c07ed0a101a4cfa54153e0498;
mem[626] = 144'h0b8aedf5010ce88e1d4b060f0d25f11bf2a2;
mem[627] = 144'h0e91f3371d6c0b6e136c09e7f17210de1351;
mem[628] = 144'h03fcfd0de78207650b23f789ed92e823e865;
mem[629] = 144'h0f88e2eef02de985042f026c1c9ef18802ae;
mem[630] = 144'h16551e69fe42fcc2e7f81627f26d0525165e;
mem[631] = 144'he09d11ece69ef541ec0bec62f8dde98e140d;
mem[632] = 144'h101ef164fbcbf7110944038ee9f91b16e3b3;
mem[633] = 144'he272f7c200d4191e014a07871a32f08af71e;
mem[634] = 144'h011c1506f4ccfa40145e1a8df30600f41e20;
mem[635] = 144'h0d3be627008fef14f6970abaf999e5211191;
mem[636] = 144'hf4411887e4ef10b4129f030dfa430614ee8a;
mem[637] = 144'hfecce3eef89711f3fdf91dd8fbb4e0f51082;
mem[638] = 144'h010d1ab4ebe906611e14fd81e3db1fd600c7;
mem[639] = 144'hefd1f931eaddf7d51df7e2701ddf112debd4;
mem[640] = 144'hf6130a4a0fb30ba41b801ae917d701bc0724;
mem[641] = 144'he7011f5ceaf011c30bcc047813fdfc4f0753;
mem[642] = 144'h171317a40d3f041ce4d50c3aeb8ee2871e53;
mem[643] = 144'h03bd0b89f3891a7f1a3be3ad00eeea800aef;
mem[644] = 144'h128512b7e00b0888e6af06aff267134d104b;
mem[645] = 144'h0226005effacf898e416edcf1294fa6c1886;
mem[646] = 144'h1610e3b607661622f61c07e80ec01cbcfd88;
mem[647] = 144'hf5b7f1dc1790ec73e555e7b0f8971fb9e5ad;
mem[648] = 144'h1bb0074006fe085e051df515ebc51150f10b;
mem[649] = 144'h0724eca81bd3f69cf93de53411a8ea6ff954;
mem[650] = 144'h026a17ba16fd1559ef3bf6f0106cf1401549;
mem[651] = 144'he6a8f272ed3df1ea1b19e36319741592fd4e;
mem[652] = 144'hf3defabbf5f71f36e5771c8e19a608daf0d3;
mem[653] = 144'h0c7f0462184b1973fc19038b1367e33af1bb;
mem[654] = 144'h025fe709166de98f0d0fe1481a24e170e73b;
mem[655] = 144'he23305b904ddfeda110b18a10c0af5400a5b;
mem[656] = 144'h1119f07f04390742f67dea49f177edeff92f;
mem[657] = 144'h1eb41be9e48f02740f03f89c0e53ff33ffb6;
mem[658] = 144'h1c1afa83141302a018d5096c016ef2fb10f0;
mem[659] = 144'he92416f2e9eb077d1a5de15d18dc0c0d1ee7;
mem[660] = 144'hf676ee01f367e06e0597f88a004bf050f647;
mem[661] = 144'h08a61ccff8d7f171f8c0f8ae09bdf18003d1;
mem[662] = 144'hef0ae1ad1b3b19a0fd3de4d60efd08521fa8;
mem[663] = 144'h0ff5e81de95be510f1b40b3ded1bf16bf5d0;
mem[664] = 144'h0d921b0a0c05fc6bfbcdf0571fabf135f35f;
mem[665] = 144'hfb4b02d7073319b1ed3af10bfad1f02e0ab6;
mem[666] = 144'hf73e09870d02fd2af717ff6e08cbe9471112;
mem[667] = 144'hf4fffcf9127ae59909bc0b7b1c0109bff07d;
mem[668] = 144'h0da4f4f01f96f37506681ce3010beffa0d7c;
mem[669] = 144'hffcffb9209e5ef53f4b90bc3187df0ac04ea;
mem[670] = 144'h04de118717b6168f17fae39601e8f46a0008;
mem[671] = 144'hec0af608e54c0eb9064f1f0cf495fe4e0257;
mem[672] = 144'hec40fec81b550dcf0313f95a0732f695fbbc;
mem[673] = 144'hf81a0c7a09aae5d0efd10de10776eefb08c6;
mem[674] = 144'h0b880a51f436e46903ff07e6f2f4039cef99;
mem[675] = 144'h159c17cc038df4a4084af28ceb28092c1bf5;
mem[676] = 144'hee17f39ef7a1edc0e759033b085bfffffcc9;
mem[677] = 144'h1d4604f7f0dff32700511a7b1e6bedc01dff;
mem[678] = 144'h00880d6deaa2fb1efd25f32f0d4ffe3ef200;
mem[679] = 144'hf20617080ce0ea79e6711f5fe6f6e9a4000d;
mem[680] = 144'h0936f0ae12df0a630b64176412ac1ca5fea2;
mem[681] = 144'h18d1f9f51fb304b20e2d067f14a70a90e8de;
mem[682] = 144'h008b19231ad81a6afd84ee6ef97af321eb18;
mem[683] = 144'h04291813173e1a32e3e61ff11a881cb61f1c;
mem[684] = 144'h0a7af224f69fe4a7fd940b310b03ffb815e8;
mem[685] = 144'h094e0956ffafe1cb0bed1d5c1a2f1f7d0a4b;
mem[686] = 144'h0380fdee0ac21174e9d80e17fac5fc92f35b;
mem[687] = 144'h0b79fc87f189046e072af20fe82d08a311ea;
mem[688] = 144'he5381ed4f98a05980420e98900af03600a2d;
mem[689] = 144'hf7b3113efacaeffa1f61fc29172800781c85;
mem[690] = 144'h1ab71224f3eb1f40ec6f1d0cfd9e1e050ba7;
mem[691] = 144'h0e6a19691295ff5ce8601b9b147c149104df;
mem[692] = 144'h14a90ed1e7b3e52feff5f8abf92a0178ecc2;
mem[693] = 144'hef8efc20f0d7e0bc178ff727e85ef2371014;
mem[694] = 144'h0ad608f1172ff0fef8571878ed67e7bff6cd;
mem[695] = 144'he03f1f5509660881190a0a0f0dc30fc3e854;
mem[696] = 144'h1b43f6721771febfec34e4dbfa29173b0e9a;
mem[697] = 144'h03b518be1d76fce4f7501d05f8a8fe94f908;
mem[698] = 144'h010a071f06e3e6320f730c9a1b3116e4e112;
mem[699] = 144'hee6d15dbe2dcf901e002e9e6ebadeddb0e23;
mem[700] = 144'h0df3f775fea4052cfe300148ed5b099ae7d5;
mem[701] = 144'h15bf12fe155a1c9bf041f46918a50e51e7fd;
mem[702] = 144'h1da9f0c6e5bc03f1f37100a7f9560a54fc64;
mem[703] = 144'h0239f4fff230091cec750c1e0e81f8d6fbce;
mem[704] = 144'he2d5165ee89dfc4af0170e9f055808dcf58a;
mem[705] = 144'h0f220265fa820d741c7f13c015d31565e0fc;
mem[706] = 144'hf06eefddf614f011ee2ceb531b370c1be8d3;
mem[707] = 144'hfab615fdfc65fa0ee3f800e6eb99f83ae522;
mem[708] = 144'he4defd6f0d90ea55fa820a960b84e1410f23;
mem[709] = 144'h083f06870cc5ef400fdb02ab01030bcf1cbd;
mem[710] = 144'he5cffdeef1600cdde3db0ef0eaf4f1d90f02;
mem[711] = 144'he1f409dfed521089175fee7ee16deaaa1dca;
mem[712] = 144'h10af1135fc71f8a619fa1760ee6105a5f962;
mem[713] = 144'hf743f4d10838fe920366ef090200ff33f44f;
mem[714] = 144'h0c32e3fef44d1ad10a7f13cf1ee516e4eb19;
mem[715] = 144'h031804dcf9bf19671c10099ae9550619f388;
mem[716] = 144'he6b211fd01cb1d0c185deaf90203e0800d1f;
mem[717] = 144'h09b0151610a4fcace832111d0ad3e00b1158;
mem[718] = 144'h10cb09c2f46b162c156e032c1ae015fe1a99;
mem[719] = 144'h15351d04e6eef6bdf98ef63a1e2ae66f0fc9;
mem[720] = 144'he10507c2e81401ecff7a1f4417d6fc22f435;
mem[721] = 144'hffa511490e7f0c3a036e1a17fedfe41be80d;
mem[722] = 144'h18ae037c0aa6f4350d2cfe65edd10df2084f;
mem[723] = 144'hf17cff0d1fc1e56b11cc1807e63ae72afa7f;
mem[724] = 144'he543f9ed1d48e5e00dcae0f1e8531822ed04;
mem[725] = 144'h0fc1edbbe3a2fd9b0fe7ebb80209fbd40f50;
mem[726] = 144'h02c103af04f10bddfb2605cb022a11430301;
mem[727] = 144'h0c41e334f88dff1cf27414fe1fdc1334fa59;
mem[728] = 144'hea1e01610e1cf8061f33158ef8fae9bd018e;
mem[729] = 144'hf7e3f7b1efad0f390930eb68e2d9f26814ee;
mem[730] = 144'h1f380e7e009307c8e6bd039b0b43e8eafc01;
mem[731] = 144'heb1c11fde6dc0f8e1b12fb2216ffe51b0dce;
mem[732] = 144'h0cd5f31817591f091079e1f9012901a4e9f9;
mem[733] = 144'hfdeb13441f56e6e5eaad08c20da2fcf7e0ed;
mem[734] = 144'h09cbfb210e6214e7f2dbe06f12f2f1fc1cca;
mem[735] = 144'hf19e1e72eb480f7ee82200ab11190d97e7f7;
mem[736] = 144'he0d9f593075a0c330034e115fc77ec27e30c;
mem[737] = 144'hed341758f8a2ee531b390fbcfe0d1aef1e35;
mem[738] = 144'h1ae2eeb1171cf33e063115eae01103c716d9;
mem[739] = 144'hf424ff44fbf105e20f7ff833e2011702eb93;
mem[740] = 144'hf3d2f01cf4a0e89617a9140ae47ffd72112a;
mem[741] = 144'h16900b0b127ae9031644f5dbe87103d3f0d7;
mem[742] = 144'hf312e607e7e811b71f6c082f0d5e100a0474;
mem[743] = 144'hf16c150412cef11de7ccf7dae4dc10e01e26;
mem[744] = 144'h1636f6ad11a11d3a1c66fde8fb930fbee7ea;
mem[745] = 144'h0259fc35fba90583103df9841f710a98e6db;
mem[746] = 144'h0f0312e01735f4fde658f08afe4ff2cbe879;
mem[747] = 144'h0cae07e01e651d54e3c7f5f4fbdd1533090a;
mem[748] = 144'he5281a62009ce5b2e34de248036713a10d53;
mem[749] = 144'hf0a3e32d073bf57fe12de1640fd6f7511424;
mem[750] = 144'hf72ff432090d11b6150906eb130906a605e0;
mem[751] = 144'h1e64f73ff955ea8df0590c8ef9b0ef00084d;
mem[752] = 144'hf7dcfd76fdf0ec4606d519d4f6aff81df49e;
mem[753] = 144'he3f70f54f4f3e9ee162507bf0c6310d1ed40;
mem[754] = 144'hf334e07110c1e2b10586ffce1a0602221996;
mem[755] = 144'h053be42ef37c1842080f189ce0a70da51fb8;
mem[756] = 144'h16c00531127fe4981430f664e2e81eb7ef71;
mem[757] = 144'h0aeff4baf2b5f80def2d167b0939ecd9e599;
mem[758] = 144'hf87014790121f95113bf10a0e011e128e4ba;
mem[759] = 144'he6511adc117807c70edf0ca3f91ce58f08c6;
mem[760] = 144'h1ecef6d3fdfdea66f4811161e4af05820a3f;
mem[761] = 144'he3fae718fac50e82fcdefb3afe6e00c81c13;
mem[762] = 144'h0d4ff0a4e080eea80a4beeb7e71617aa12e8;
mem[763] = 144'h139ff5eef4711487fcc61fd61e590f40152d;
mem[764] = 144'h1909f0541c93f62008e118a5e8edf2f6e26e;
mem[765] = 144'h1294eddfe8eb10b9e827e5dbf04b02b70623;
mem[766] = 144'hf0afe709f694ee6c18e91b52f046f44df5b7;
mem[767] = 144'h0253eda3f67d1993ee25f58518a61c46f32c;
mem[768] = 144'h1198f4df03e40bf4f47ff5f1f19bf9bdf13d;
mem[769] = 144'h011c1abd04bc09c5e3bde9ac1081ed8b11e7;
mem[770] = 144'he4b21111180e01c91dfc10cb0b86180cf64c;
mem[771] = 144'h0c1efd3fefc703690eaa023a1deb04cd014e;
mem[772] = 144'hfe5b13bc0afaf135eee00dcb037404720747;
mem[773] = 144'h1e00089615b9fcf8f59a1db8fa1107090be6;
mem[774] = 144'h022bf7fce52de19c032eefd5ec39164de554;
mem[775] = 144'hf86ae57d120815c2ef750947f5401ee6fd7b;
mem[776] = 144'hff28115407c1fe98e50010a813b21065fb2e;
mem[777] = 144'h06a201f41a17f91ce154067e1b6c0807fa66;
mem[778] = 144'h080ffa720598fee80b96f0c41e2c02690e64;
mem[779] = 144'he9a2e3950adff46bfce7ffec15d2f719169d;
mem[780] = 144'h0c6904d51c76ff49128beedf187ee5451981;
mem[781] = 144'he8eeeab409d5f86aedd611dbff78e2d71eec;
mem[782] = 144'h1d70e8c4fff5094fe8db09c10db2e9e91331;
mem[783] = 144'he2aa0686f384ee61f9cffb380f20f1191bb6;
mem[784] = 144'hf5b1f19104d812ebfc9d171aebf4f1080523;
mem[785] = 144'h0b47e372ffce0f4202b9ec07e200106c16dc;
mem[786] = 144'h111de16617c2f063053beb8300f5f929ff20;
mem[787] = 144'h174a061e1d7ef32becfe192018d60f6f18a8;
mem[788] = 144'hf4c0e33ae704e290f62a1d5f190317f5f621;
mem[789] = 144'he02ff6c2ff0401b81db402590c45127a13df;
mem[790] = 144'hfb4c1a62f7b31d6913a2ee250f1b19c0eca4;
mem[791] = 144'h08891b4700a1ecb0e46ee19f09d50b15f01a;
mem[792] = 144'h1bb0e6c00bfd1dd6e0d6eb0de577e40a16e3;
mem[793] = 144'he716e8e9e81e18b7ec94e5dc0b9dfe9011d3;
mem[794] = 144'hfc771c271653e60c0ab607a5fdbfec93e5ae;
mem[795] = 144'h0c261138010fe8520775127cf93bea6b0e98;
mem[796] = 144'hfbefe5ad0cec1952e563e31ae7e50cb9ef2f;
mem[797] = 144'h10d7f54a0ea405db08efe1d71d0f1cf4edbd;
mem[798] = 144'h0f63e93b0f0fe3ea0ce90bbdf82e13da0087;
mem[799] = 144'hec1c19e5e096143201290adbf8da1bd50cc7;
mem[800] = 144'h0e45ffa3e783e0ee031f1d6d19970ee8ef5d;
mem[801] = 144'h03931b69e9b3003cf914fd15ea651f69ec15;
mem[802] = 144'he570f929eb0ffa28e6630c44016afd510b7d;
mem[803] = 144'hed7fe70cee43196812e1e694e32e103c097d;
mem[804] = 144'hfd71e9850e550f9f1d7b007a057eef750e40;
mem[805] = 144'he51ee9c4eef1034ae92f18cf0c7fe3eee9a6;
mem[806] = 144'heeda15b80b17fe1afd27f2041fb70b421920;
mem[807] = 144'hf5d318d3f072125ef6b0f30eff92f252eb64;
mem[808] = 144'h0217e51bea9f1b5d0dc81dae194ffa761d4d;
mem[809] = 144'hebc3097f1f021d74f09d1cf3fd20f557fbc8;
mem[810] = 144'hfb61f6e8e9a51af2fd96e5b60ab915ffe4a5;
mem[811] = 144'h0c6df8331f3c11bcec89f795f03516f3f949;
mem[812] = 144'h0a0c011cecb0fdc81c8fe9c1ea9d10f202f8;
mem[813] = 144'h11080c92fd4c0054fc19e767f9010952fc02;
mem[814] = 144'hea220c5e01331976e9f6ff7d07faee57eeed;
mem[815] = 144'h0d9d16d412c2073719bd04a8152304e2fabd;
mem[816] = 144'hf008f187fa5ffe7302b003d60a26f3c0e08a;
mem[817] = 144'hf92c18f0f111e5b40af30eba0b2509b5fb90;
mem[818] = 144'h0ea4f02a166a1ca4eaaa1a86e696ed540d10;
mem[819] = 144'h006ff601f95212d61e5fed920ae50387fdd7;
mem[820] = 144'h0b26ff73187d1c78f3490aa30205e786e781;
mem[821] = 144'h0455e568ee1df546e6a00ffbf3501f4cf416;
mem[822] = 144'he1d205f2e1b018a0059511c3ec9ee2990b1b;
mem[823] = 144'h0861ef8806640275fb1319f6e17ef13e05b3;
mem[824] = 144'h0cca1d54f148e0db199a185c184918f5efa6;
mem[825] = 144'h007e1d49ee5a04fe010bec01e5eb192fec1a;
mem[826] = 144'hff3be414f578f9a51c8af415e297f495e149;
mem[827] = 144'hfb03e681ef901c0b14b011e7fca9e202e454;
mem[828] = 144'h1cae1d65e0bb1b711231f6f4faa8e4411333;
mem[829] = 144'he569fb4cf05c12acf0b6e465f332f994fda0;
mem[830] = 144'hef24084c13c7f2a3e69ce1a1f570e6591053;
mem[831] = 144'h0b90e53b05f3f8c2f4cfe6e70f261481f47e;
mem[832] = 144'h053d1692fb581f4ff00ee887fbedfeb9e801;
mem[833] = 144'h0149fa1ceee7f8a71e61134bf539f8cbf031;
mem[834] = 144'hfcaaed121d6a1ad6e689ea691fcd1077fd7f;
mem[835] = 144'hfb34f0e6ee5f11a7fae40ce71e811342e619;
mem[836] = 144'h04bd1912e008ee2be9defb7c0938e9b1eb92;
mem[837] = 144'hf5980f48f41dedc21a27e8f2154107c7ff2b;
mem[838] = 144'he1aae62409b717851fecfac2eee8ffb506df;
mem[839] = 144'h09cdf99704220094ffc50a20e29b0066ea36;
mem[840] = 144'h0bcd1a230044e146085c067ee70018131074;
mem[841] = 144'h00400a830e4bf4c8efea1e431eb6f71be514;
mem[842] = 144'hfca21174ed4ffc690832f1a7089518a5fd90;
mem[843] = 144'hf326077810bfe06304c9ec1afa00ff5bea92;
mem[844] = 144'h1159ec9b1ae6e1a7ee840f24ffe71d2f19be;
mem[845] = 144'heccc068218250c761714f7d812b8ff8bf88c;
mem[846] = 144'h01661d89067101611d49e464011213bf1c89;
mem[847] = 144'h1231edcdfb63fa2ffaa411e009a70956efc3;
mem[848] = 144'h1b50f24fe88dfcdd161e04cae2afe6cbffd9;
mem[849] = 144'he1101849ff1e0a73edcae1c0fbb1f949fa56;
mem[850] = 144'h09ae0a63114be7c2e95cfb66f6f902fdf750;
mem[851] = 144'hef570522f1480655efbaf720ee190ae71df1;
mem[852] = 144'h15f1f409e68606700fa5165efa15e3cfec68;
mem[853] = 144'h06d915981fb5e98be75fe04b114f1e5c0d08;
mem[854] = 144'hf18eef41192117200ef1e6eff5740bf0e34c;
mem[855] = 144'h1aabe6acf6af03a50e5ef354f9da049df9b5;
mem[856] = 144'h1d90f7b7ed2ffbf9f156e163e4a51c271e21;
mem[857] = 144'hfa2212ee16dbe2b408c7f716f29d02d01a3d;
mem[858] = 144'h07a5ebe40068e44be187fe4b0d7702bce810;
mem[859] = 144'he953efd80a5a1b0706bdf3151948ede31f37;
mem[860] = 144'h188916c5ffcee400f81114df15de074617bf;
mem[861] = 144'hf39b1d5e0c3d0f74e472e7ceec2b0567f8f8;
mem[862] = 144'hea36069ce13a0627e0c0109e16a1e15d12cd;
mem[863] = 144'he144e5e209791e650d4efc3ef061ec65eda6;
mem[864] = 144'h0329ece6e3cb0945ff2eff11eaa8eb380d74;
mem[865] = 144'hffac11de0786054ff1adf14508901a030efe;
mem[866] = 144'head91a8b180005e30afbe2ae0804f6dff1f0;
mem[867] = 144'h107bfbddfac803b0febce017e561023f07b0;
mem[868] = 144'he4daf21af7b4fbe9f21b09dff0baecd0f713;
mem[869] = 144'he7f7f785ec1b03df0fac12a41f2916b30655;
mem[870] = 144'h0c72e17ffd25f8cffe5ffa8de8e6e27700ee;
mem[871] = 144'h0dff1d37ea4ff46b1b00052cfe0cec4908e5;
mem[872] = 144'h0dbbe63ffcf6e35eec33eba3fc03f5930c2e;
mem[873] = 144'h087efb20f29cf9610c7c1ea4f45debcff77e;
mem[874] = 144'h17461a5713c60278e123e433ffaffe421004;
mem[875] = 144'hfe321edce28c1a0fe9d70766f043f0deef96;
mem[876] = 144'hf5f303c5ef38ec1a17070a661c92fedf0646;
mem[877] = 144'h0292fc74f26f1d83021de2b0eb720e2bf12d;
mem[878] = 144'h16ce1141f037eb4feda1e300028c0f880fea;
mem[879] = 144'hfc00ff781940f319165aeb29f547efa5014f;
mem[880] = 144'h161302b3089a12fd138de16707e60c390eaa;
mem[881] = 144'h1c111dcefbc10e741e85fe0ce04d05b80a99;
mem[882] = 144'h0203e071e451f70508f3ee73f92d0cdde4e1;
mem[883] = 144'h12affa911fdaf32e0ad1f899f6f80be6e9fc;
mem[884] = 144'hf0a1e4241a8aeb1cf50c004606fd1791f9e2;
mem[885] = 144'h0539e822166ef5080e6100e5072ee284e367;
mem[886] = 144'hf51fe9d71750f7d107661a62f58aeffff2f8;
mem[887] = 144'he73aeb31017efa530c3ff7b91d0b05e80cd0;
mem[888] = 144'h0f7df788137916d11ee5f32018e5e5f20629;
mem[889] = 144'h108be9621d710ebb10aee904061f1db91824;
mem[890] = 144'h0a720151e1720374e3671200101de563093b;
mem[891] = 144'hf3511a4be033f3ddfb94eeb5f003e36c1ba3;
mem[892] = 144'hf403fe0dee5ce86110300d7710ace1c1f413;
mem[893] = 144'h1a3ef0770c850511195105cbecd60bddfc93;
mem[894] = 144'h0e02f926e5851490ea8f08841aa5fc9017f2;
mem[895] = 144'h145fe239f048e061ecd4042b01c4ead309b8;
mem[896] = 144'h18f2ed1712ae0af5f84cfdae0de6e19f11cd;
mem[897] = 144'hf23a0058169af33ef1aaf4ecffce1b61e087;
mem[898] = 144'h08900fc509640e09f7d60aa2e07ee6fdfc75;
mem[899] = 144'hf8b2e3781a4c030a168af47c0eec1d22f97f;
mem[900] = 144'h0c01e3df1fefec79e016f79608801156ee73;
mem[901] = 144'h178de4b1160209d6e7d2eec7f767fc821e24;
mem[902] = 144'h100818560ffa0743e82b0414043cf43def4f;
mem[903] = 144'h0bd70096e9e919e212f7ead2f27efbb6fca8;
mem[904] = 144'hf2100c2f0b0d14a4fa4202c50510ffbffe38;
mem[905] = 144'h092dfeeaf8f206d8f0b4f02d1a3016e4018f;
mem[906] = 144'h0a810e221dc1f0ad1133f212f6c0e6b413c9;
mem[907] = 144'h085cfd95e861fed8f4defff10cc3e0fae6ac;
mem[908] = 144'h007e00181166eb2af5f6f21f041b10dfe303;
mem[909] = 144'hf76afa32046f1daf03821ec9069b1309fa6e;
mem[910] = 144'h065b0f7ef032f80d18d41a4f17ee110205da;
mem[911] = 144'hfa68fbf6f931f71916421b66f1671456e438;
mem[912] = 144'h1979e0b7e5e2f8e0ebb601cce0d6e4d2177c;
mem[913] = 144'h0ce0fb08e97e1e7efef91e35f8bbeede0d0d;
mem[914] = 144'he0e7132ef4b90172ea6b17c402e6e06cea9a;
mem[915] = 144'hf45bf09e03301f5d1c60f9250689082d1879;
mem[916] = 144'hfbae050feae9ec1a04170bdb10981ba20ad1;
mem[917] = 144'he85d191a01d012a31eeb0ce9e9a6f4af04b3;
mem[918] = 144'h12ece795fc6d09ba18891293fd80ea9c112f;
mem[919] = 144'hef36fb0e19ec17721595e2a70a21e822f19d;
mem[920] = 144'h17b11a9df0e0feaf07ba0d271e35e5ece7c4;
mem[921] = 144'h0f7f151c07270dfdec5beb94f739ed88fad4;
mem[922] = 144'h083f1a6af61e1a0905911bd8044b15edffad;
mem[923] = 144'he37ee631faf8053d0d04069dfec6103b1cb9;
mem[924] = 144'h00cd1679fa9bf830136102d0043a1b72fa26;
mem[925] = 144'h1501151f19b61f9517b21b60e9d8f2ee0601;
mem[926] = 144'hf8191db2107ff6b7f2e00d7afd3015c3017e;
mem[927] = 144'h01f7fde60279116dfd721cccf6a514b8efa3;
mem[928] = 144'h0239f826fad804e5015700ee0c71052c1412;
mem[929] = 144'hfb67090c1bf0e01d11a4e3bf0237fbcdef28;
mem[930] = 144'hfe1a1a1908fbf0b1f8eef6100095063af985;
mem[931] = 144'hfec7efa00622fee9e83aeb99fce3146c027f;
mem[932] = 144'hf4b81591eb0c1b83fc6de659eef8e52b1d43;
mem[933] = 144'hf747ef070a8d13e3ed4e09a41e72e9d904a7;
mem[934] = 144'he37016e60656f265ea9df3bb190efd6a18d3;
mem[935] = 144'h1835089a0cd81b0be3031edf0aafea1be3f8;
mem[936] = 144'he7da03eee11d09c01b3be23b0498178dfdcb;
mem[937] = 144'hf76af3a611e1f01d15c5fa55f1aa00eb18d6;
mem[938] = 144'he57a1b46056be0acfa971a9d001318c51edb;
mem[939] = 144'he0ef13c81ed5efc61c8ee14fe6b707cee19d;
mem[940] = 144'h053ce6341152fd3b062e0dc6ff2cea5ae804;
mem[941] = 144'hf11200c5e519f142fe69f0a4160b1221fd98;
mem[942] = 144'h01c8f7b2fc09fe801a6313d9fb2f0a4ceb62;
mem[943] = 144'h0c2f1f1018bdfc89e586f2410ce804801446;
mem[944] = 144'h141e15c6ebb3e0a0eb3a19821974f95aedf9;
mem[945] = 144'h011f1a3ef58a1deaf28ae07d0c7cffad0935;
mem[946] = 144'h18ba1e5f184eff8f1333e1beefcb0a301aea;
mem[947] = 144'hf1d30d62e50a0bcb0c8eed651a6bec1802c6;
mem[948] = 144'he2f3f63ce699ff65ea54e30df27ae479fba0;
mem[949] = 144'he5b3111af7a80bb5effd178e0d3317ef04e7;
mem[950] = 144'he097175c0cb3e677ee1fe618e7831a8ae2ee;
mem[951] = 144'h084b02ff1bc5041416d0056fe0a3ede20139;
mem[952] = 144'hf90d05cd07f7f05d0872f76df42ee6c30bba;
mem[953] = 144'hf976199ef3d7e36aed9fff3e0000e346f84a;
mem[954] = 144'hffa7f806f2bf0e5a143e04d311aaff1df91d;
mem[955] = 144'h1a5700ed1788fbaffe65f139feda02130c2e;
mem[956] = 144'hf3610f49efe90eb1e68f1b18f8271babeb9d;
mem[957] = 144'h1d861b53e9bb04f60df6eec00496f2e0e239;
mem[958] = 144'hf268e03b02fae2a01f5c1dd6fc110515fecc;
mem[959] = 144'h07b71e7bf03006581daeee721d9ff9c21efe;
mem[960] = 144'h16dc0c651f9af822e4bee9b60da8fa24f014;
mem[961] = 144'h0d03f4eb0122e9db1687e5b3123cf786f6bc;
mem[962] = 144'he74ce7acf7e916c6f99619f0e2e8051f00ba;
mem[963] = 144'hea1d0a2a04e7feb8e51f05ffe0341018fc51;
mem[964] = 144'hf3ddf64d06cb12f70d0617a3e1741e8c1372;
mem[965] = 144'hebb2ff2cf451f215ff1ef6421110f6890674;
mem[966] = 144'h0e99194eeeebe1510833e512e6cbe31f0393;
mem[967] = 144'he39ee84301aeebedf9cb078f0dd4f2d10394;
mem[968] = 144'h1171f65e0b120b44e9d504a6139d08f2fac9;
mem[969] = 144'h04a202531e3410940e1b12cb02d7fa80f770;
mem[970] = 144'hf99906abe82f16d014791ec309fbfefdffed;
mem[971] = 144'hf3bd13a303e706f001f50cc516a214b7f0d4;
mem[972] = 144'hef68eace131315d10f33069de535f23f148d;
mem[973] = 144'h194009f31045e5f902e81bca0fb71c0be9c5;
mem[974] = 144'h17a7e5c11381fcabe285fb57f08d05f8f62b;
mem[975] = 144'hfeb9efea128ee0fbeccc02bb0ef7e4d2e8e3;
mem[976] = 144'h012ce031f0ae12fc1e83167ff69d0d9aff95;
mem[977] = 144'h0163f5d51e0706111c87124ce3f309a7fb99;
mem[978] = 144'hfc53013711120e5d1054fe2615df1a3d1a81;
mem[979] = 144'hf94ee7a1197c0fc7e6a1060c00a5ee2eebc3;
mem[980] = 144'hfb4ee2a8fa5cebd402d109b8f2a701641316;
mem[981] = 144'h073712f913dc0153f2bcf529eb5af996e8b5;
mem[982] = 144'h0a85e0c0fd10e988ffa503cbf915f20be9ba;
mem[983] = 144'h0cc7ffb1f1950b4d040bf1ecfe3111f513c2;
mem[984] = 144'h1563f46af9a9f109eed5f581fe92f58bf674;
mem[985] = 144'he5b7e446140f124d064104cf1fbbf57aedfd;
mem[986] = 144'hf0fb068ee01c017afc72f0b91089e3aaf7ad;
mem[987] = 144'hfc93e1ac09b1fe75ebc7fee2fd66f07ded26;
mem[988] = 144'h0ddaeb5efdcfe8d2e0d4fac4061cf01ae035;
mem[989] = 144'h1ab1eae40900e68cefbf1a7607c0e7bbfe86;
mem[990] = 144'h00d3e7430274f013f14712cce0d7f4c00af5;
mem[991] = 144'h042906bb1b3f0e5ff46ef2a5ee2b156b0b2a;
mem[992] = 144'h0c83f171fbc9f085ef97ecc5ea9de229ee7e;
mem[993] = 144'h048f1ecef523e7cf061fe96819d3ede014e8;
mem[994] = 144'h0a36149beac1ecbcf2e41a45e31608b4e5e2;
mem[995] = 144'hf245e844fda3ed7ce85eeb08e93ffaa7eff3;
mem[996] = 144'h0765f90bf05eee94f04c0712f6a912691fb2;
mem[997] = 144'h1b4df3c0e691034f0dd1f2caef651a4fe23c;
mem[998] = 144'h057612ede2ebf504fd5af6f50c9614251f20;
mem[999] = 144'hfb8d0006eec2f6dee0d019bee5a3f4b706cc;
mem[1000] = 144'h0089e0f918a416fa1c0ff0190812f429eccb;
mem[1001] = 144'h1530eb1f1cdce561e983fe6c0d70f62218b1;
mem[1002] = 144'h19eef322eb9805de1ecaf82412aee3e3f03f;
mem[1003] = 144'hf91209eefae4fe661dff01bd1dd012fb1a4a;
mem[1004] = 144'h1146f51ee6da1d021bc5e39004b2efdbe318;
mem[1005] = 144'h0f99fae11e2a1044123a1fdf149416de104b;
mem[1006] = 144'he7c7e07b1e85f0cce12313661b5dee7504b2;
mem[1007] = 144'hfa8e1336f5e0f0ca0f42143b187aeb3af848;
mem[1008] = 144'hfc6ef72413fa18cdeff6f69d17afeb61f091;
mem[1009] = 144'hff5f07021fe6e06a0a82f6dc067e1563ea6f;
mem[1010] = 144'hf2de08c50143ea1108f6f4fef43f01a31f8e;
mem[1011] = 144'hef8ee4fdf97fefe700f71bb6004c129ef23f;
mem[1012] = 144'hef8e1772ece81663f929fb010994f3d3ed8e;
mem[1013] = 144'h0f3f008ded9efed304c0e0da19e3f97cfa7c;
mem[1014] = 144'h1ad2eba8071de218e68d138a18de1929019c;
mem[1015] = 144'hef04fb5df3f1eb881244fc29fd19048d0077;
mem[1016] = 144'h1fe4fa99fedffbf4ff850418ed8c16a1ec80;
mem[1017] = 144'he422e450fb07110904ac02701132e326f974;
mem[1018] = 144'h1347f858f156ffbc04201212e10cec5bf3db;
mem[1019] = 144'hef48f65fe990150603981ca6f0190cadf291;
mem[1020] = 144'h12a4edbb167c0b87eea91d1cecd0ebe4114f;
mem[1021] = 144'h14cee7210f14eafbff090a9806b90db1e13f;
mem[1022] = 144'he8beecdbed32fc17ee61e0830f7af66b0726;
mem[1023] = 144'hed92efbded7bf155e1e70f8aec09feb7edc7;
mem[1024] = 144'h1cd4fb1ffa92f17a1527e2bae9d91a12ef39;
mem[1025] = 144'hf74218e3e188ed56f139f5450d92e8c8f58b;
mem[1026] = 144'h1cd31d0d0829f7ba18a60c3b1224f09ee62c;
mem[1027] = 144'h091f0f0fe6b2e64afedde39b045ef99901e5;
mem[1028] = 144'h1610e19eec04ffa3efa8003d06e3e796f50f;
mem[1029] = 144'he05613a8fc92e9200d94f1e90ef7fe66f173;
mem[1030] = 144'heab6e20ee1130f04e5cee2ffe2f51286020a;
mem[1031] = 144'h0a7a06a4f767fa76ff13ef88f7a707f502b3;
mem[1032] = 144'h0a831b81fec81991ff1713a0e2b10467ed5c;
mem[1033] = 144'h05c41499f7b011f1f9d1e2960d47eecbe915;
mem[1034] = 144'he86bf21de7e9e3ec1c141e4c0e91f6cc13b8;
mem[1035] = 144'h1a5b1964118cf7ac1f8b07fe1dc8e0aef113;
mem[1036] = 144'h0eb9e11603bd0281099bf78207d6146bf352;
mem[1037] = 144'hfd43e4d0e39bec0000c703990dbc118812fd;
mem[1038] = 144'h11811b261b240ead1658fee90035f6bdeffd;
mem[1039] = 144'he6b4fcd6f84808280b7c1e95180d0a5d0830;
mem[1040] = 144'hf66b0d6afd16e0df1684e99e145f05bfe550;
mem[1041] = 144'h1e07f69515a001e8e2f012b0e8a6e4a21082;
mem[1042] = 144'h0c6f1c9a0db0172ded69e11e1e3ce346f40a;
mem[1043] = 144'h1d3e039709bb0d55fc82ece70919e2e303d5;
mem[1044] = 144'h1880eaf7188f1f16054bea811065ff1110ca;
mem[1045] = 144'hfd061005f8bdf5e0e66016e217fb19390c21;
mem[1046] = 144'h1e34ea6f07f4fc3a19cb0828f2b3e1940df3;
mem[1047] = 144'h05d9e59b1fa71343f53de2c81c86f596fcff;
mem[1048] = 144'he61bf55c1a271aa2022b1b93e5dcfecde786;
mem[1049] = 144'h034ef20609d212a8f593fd840e17ed851435;
mem[1050] = 144'heb81fdc70f4308eaf3730a47082c1bc2f4d6;
mem[1051] = 144'h0d63167b0e12115ef8b6194400d11cd70063;
mem[1052] = 144'he31a0acd18661c0b08a9e791f555024007b3;
mem[1053] = 144'h0973fd7505e2eb581be7166c1d74e599f109;
mem[1054] = 144'h1d98ed2ee6aaf9fa0468e114e1a1e677084d;
mem[1055] = 144'hfc3cf70af230045f168103b2ed39e4e6f52d;
mem[1056] = 144'h1eebf858f86bf928e244eebe0985fbb2e744;
mem[1057] = 144'h1326f7df189cfb6c17a515970734e7420e24;
mem[1058] = 144'hed3c1dddf39c0bd4febe00ca05890ed81244;
mem[1059] = 144'hebed15661f7716c513170087ed3eecdefa92;
mem[1060] = 144'h1b69152e0869eb06e360e5f71899fa94106f;
mem[1061] = 144'h036317271194175bf417e9adf1230c001f0c;
mem[1062] = 144'hee0e0301ec18f9a4f989f5b31d0ae50c13fe;
mem[1063] = 144'h105bedc9e9caf015018de7cdefbc1fcff11c;
mem[1064] = 144'h0c79f35cf4181945197a156f069f08a80805;
mem[1065] = 144'h1a2c1364186d142003290dec0d82ecfdfd5f;
mem[1066] = 144'he031f29213c4f4861626e5e0153f0502ff78;
mem[1067] = 144'he85ee95fedf2efb1e0d818ed1967f97f052c;
mem[1068] = 144'hf253ff6cea5efaf607f30ac0f5870ad1e7b1;
mem[1069] = 144'hf681e424177f0496f82d0e990f4bf87efc5e;
mem[1070] = 144'h0a48ffe1e851ee05ea170f3e1087f901001f;
mem[1071] = 144'h0977168d0b7ae8aaec511f4f010df3570b1e;
mem[1072] = 144'h04821977110b022dfcad13ac09dae7881a71;
mem[1073] = 144'hea40fcaafea315b4ef7b0af6132703b0e2a6;
mem[1074] = 144'h0381e44ff0e00897e73bf53c11cbea84068e;
mem[1075] = 144'h1a36e6cb0b66128001da1097f5c6e2be19f7;
mem[1076] = 144'h0402e0d207d61cce068c0bdc19501a9d1d86;
mem[1077] = 144'hf7150369fe5aefcb1b69035c16840a3defcd;
mem[1078] = 144'he273112d005fe5eae191e06710b41af017f1;
mem[1079] = 144'hf4edf73115460a8f12f7ffd512c70db71511;
mem[1080] = 144'h06e2e8c4f1d1012bfeeb19fd08aaf0531da3;
mem[1081] = 144'hedc7e807142f05e416c7063b16af0cedf096;
mem[1082] = 144'h1c9c150f022c1f8f008911f5ea7ee3911dd7;
mem[1083] = 144'h0f5df01dfca41329fbee013511a4e28de1de;
mem[1084] = 144'h0980faa51ab60893eae8ecb0f930e952179b;
mem[1085] = 144'he26907ccfa250312e9f4ef7ef8d0fed7ec14;
mem[1086] = 144'hfabdfea007e3f792ecddf2b9f3b8e7f70571;
mem[1087] = 144'h06ed194fe8781905e27dfb5ee971eb19e241;
mem[1088] = 144'hf6fb087df049eab3e5fffea0f5f80d9fea0b;
mem[1089] = 144'he8f1fd5010950f610a7502b113a3f32de9b5;
mem[1090] = 144'hec03140408dd1a2d13c8f257ee8705a7e1c0;
mem[1091] = 144'h02cf1d19f4c6ee842033fbc7edee221618ce;
mem[1092] = 144'hf3edf9330b9de6951cebf3300c6fe1efe265;
mem[1093] = 144'he656eb27fe800cd5fb880c23ff53ea59ee1a;
mem[1094] = 144'hf94117b30afa19fb23e1028ae773f108fa05;
mem[1095] = 144'h09ab05bbfa450943f60af1040ee8f2240621;
mem[1096] = 144'hfa01f744111c1cbde96c14e4e96ffa41fcfd;
mem[1097] = 144'hf5d9f4cefc3f0028f224ea1f1aabf2d2e94c;
mem[1098] = 144'hf171f6c11c58f2bd1e3913541246e4730c99;
mem[1099] = 144'hf338fc4fe9491950024deaede881ed73f133;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule