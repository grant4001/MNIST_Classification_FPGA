`timescale 1ns/1ns

module wt_mem4 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h05bef09408a4f994fdf90a010e00fc71f6c7;
mem[1] = 144'h0702f312f4be08a3f75e0a02fefa0d4200ee;
mem[2] = 144'h0163f5e5fbaaf95905db03ea07a3f5c208c0;
mem[3] = 144'h008803d1fbb0f744059c0f84ff7dfc6bf0f8;
mem[4] = 144'hf1b6fd27f935fc8b04f0fdad00a103ecf053;
mem[5] = 144'hfd61f57f02f8f9d9fd57fed9f4f3f2d50616;
mem[6] = 144'hf7890842f2c70d24f5cd0245f86df8fa05a4;
mem[7] = 144'hfae6f821f788f48ff129fdee028007e005c3;
mem[8] = 144'h00b9f7130231ff24ffc00add096e0cbd078a;
mem[9] = 144'h0f58003ff4210b4df58cf0e208f5fc960dd2;
mem[10] = 144'hf9840846f26bf17a042208b1002bf2d70cf6;
mem[11] = 144'hf753f4dbf96604890904f798ff7ff33800fc;
mem[12] = 144'h0f90fc78fca5f54cf2220f38f81905b9fca4;
mem[13] = 144'h04b30d40fde30d9f093ff813f505024907e9;
mem[14] = 144'h09a5010a0f810f61f2a4f202f0be09780de1;
mem[15] = 144'hf5a90ddaf3170a72f360ff9f084df5a2f608;
mem[16] = 144'hfe5c0b39f42ef7adf8cf0a8d06ca0734f451;
mem[17] = 144'hffdcf42708fd047fff0008d5f9c0fb8e0565;
mem[18] = 144'hf8d9fc440aa30c73ffce037d0a4506290255;
mem[19] = 144'hf6420eca0700fe6303b8faf5fd8b0602004c;
mem[20] = 144'hf54bfdf5fe730dcd0df20acc02ad04d600de;
mem[21] = 144'h0b43036302d9fcb00cf3fa71f9f90ce60b1e;
mem[22] = 144'h0740f3b1f912fbecf1c402fa02830f3a0ea3;
mem[23] = 144'h06cc0b43f829f9f80d26f2c9f95304700ac0;
mem[24] = 144'h00700ea30dc90f990593ff4a0b1efcd9f765;
mem[25] = 144'hf0c4f3dcfb3cf687f02008e2fe850733fde0;
mem[26] = 144'h098fffba0a66f1f40800f4da0e4b0793fe73;
mem[27] = 144'h07a60a4a0c2a013a0184fb13faa00e740142;
mem[28] = 144'h09740abe0213f344fb28062f0a31fd870784;
mem[29] = 144'h0e8205fa0c27010d005dfa46f0baf19df716;
mem[30] = 144'h029d0bac00b90466f1cb060304d90a1ff697;
mem[31] = 144'h0d770cd202a6f47a00090649fabd03bdf0ec;
mem[32] = 144'h0978f3990d74f7770081ffee033a0acff8db;
mem[33] = 144'hfc74fab60a96f2c00af3f5bc077cfbe8f42a;
mem[34] = 144'h028200e9083ef556f7fd0c5307200d26f21f;
mem[35] = 144'hf44904a1f070fc7d0c9703e40f32ff49f75a;
mem[36] = 144'h0669080504430a620e66fac4f0e3fac2f6b7;
mem[37] = 144'hfee00501fe0e01080c3df8d4f1acf3430f4f;
mem[38] = 144'h0c8901f7f118fb2a0bc1f44ff3bffae9f24c;
mem[39] = 144'hfef20e200f6effc90f31fe5ef9d60058fd8d;
mem[40] = 144'h0cf701f505cb04500d9bfeb6f50008dbf840;
mem[41] = 144'hfbac004cfc7e03b00f6c06130fb5f710f1ff;
mem[42] = 144'h02f4f833045afd9cf2ddf40a072ffe3ffe52;
mem[43] = 144'hf3a0032e05e0f12d00620e11030bf0220bd1;
mem[44] = 144'h0a320d690e17fe5f079e0042fc2107910950;
mem[45] = 144'h0764f7750ab2081800a8050cfd0ef7020a10;
mem[46] = 144'hf65bff520bd5fa94f820f1a8021c0248fdd1;
mem[47] = 144'hf2f3f484fe160e5ff4a60506f495f28e0a3b;
mem[48] = 144'h0b8a08d3fc3df8f50e56f50203730d30094d;
mem[49] = 144'hf2db0217fcd3fc0d0eff0faeffb5ff7ff818;
mem[50] = 144'hf505f3a8f31109ec0bf90cf1ff3c0437f0f4;
mem[51] = 144'h062e04460b990ec20236f56401810d9af5b2;
mem[52] = 144'hf3bc0c0bf2070d6efd670d5a02d1034d0467;
mem[53] = 144'hfdc90a1defd70240f3d60e380202f98e0876;
mem[54] = 144'h0a720c29f8880dacfc3d0b95f550fc0c078e;
mem[55] = 144'hf1150f8e06f7fee4fd7e0273f49d0e630121;
mem[56] = 144'h0ea602c7f92ff2a80cf4f16b096ff300ffe5;
mem[57] = 144'h0233fdd107fa0ac5f495093fffd4f0c2f959;
mem[58] = 144'hefcb0bb0f8dbf48d0301fdaff887fa0a0cac;
mem[59] = 144'hff9ff93cf1f5f512019bf513fa30f1e60e06;
mem[60] = 144'h010ef2d50035ff380bf605930959f0020209;
mem[61] = 144'hfcc00e3a0c1c0e33faf3f6b90d00f93df438;
mem[62] = 144'h0f5309a1f4080c9801b504e60bb0fd670b9a;
mem[63] = 144'h08d607fe0f1f07320ad8f36a0877089afc9c;
mem[64] = 144'h0ca5f4d50100019cf7ebfb58fda9fe5008be;
mem[65] = 144'hf751f9b60e47f79e0a60fc8c04500c36099f;
mem[66] = 144'h0f070ba7006cf92f0ac903400912f433f15b;
mem[67] = 144'h0411048fff7f06fb043df99bfbf3f209f1f6;
mem[68] = 144'hfe49ffce09050f300c1c038c001af1e90d87;
mem[69] = 144'hfa25f0bf0744f982fefcfa04fb7dff56f0a9;
mem[70] = 144'h04ddfa3af891095ef68108d5fe210318019c;
mem[71] = 144'hf4d40c41f1b3097a0c6908ec095b0b34fdee;
mem[72] = 144'h056c032cf2ed0df0fb25f58cf151f1e3f738;
mem[73] = 144'hffb9f54df37a0ddc07ae0101f363f9c90936;
mem[74] = 144'h0a15f8e503a9f2cbf76a0e57f0caf96d0801;
mem[75] = 144'hf2dcf838041e080202bc010006ba0e910af5;
mem[76] = 144'hf5f0f72df110f7fff3320f22f73a007cfe2d;
mem[77] = 144'h0190f33100650b2a01810dd7029108f1078e;
mem[78] = 144'hf038f9c9f086f202f6e40c1df3d107d1ff5e;
mem[79] = 144'h0aa90b05fef90a97f36afd3908d0f01102a9;
mem[80] = 144'h0524ff1605d602b4004f01ce0315f36c09b5;
mem[81] = 144'hf3f001e3f93afc7af588f113f6d3f6fe063d;
mem[82] = 144'hf312fdeefc660d940885036ffddff158f8f2;
mem[83] = 144'hf6970927007d0890f4b202a7f84d05b205ff;
mem[84] = 144'h0edc00fef54b0d81003affafff510889f858;
mem[85] = 144'h0608f7500522f8b002370273f47e07060a85;
mem[86] = 144'h0879f2d4f020f9bd04f1f016f6f403d6f790;
mem[87] = 144'hfd86060cf967fc67f19c0f0c0014f0e3fbb2;
mem[88] = 144'h0927f1fef6e6f99509e50025ff3605f7f6cb;
mem[89] = 144'h0ff9f4b7ff33f510f4a30bb80294f7b0f95e;
mem[90] = 144'hf1f9061ff466f024f85af4bffba2f76e01ed;
mem[91] = 144'h0cedf16c0271fba20bdefe240ae3f0d80cde;
mem[92] = 144'h0e5f09f7f6770346feb9f6750477f5d10647;
mem[93] = 144'h0bfafcec0d8df1290524faf70683f521f470;
mem[94] = 144'h0e250c12f6080f94f9870f44fd56fd01f1ed;
mem[95] = 144'h0777f9b0f5caf0ca02730510f527f750f7bf;
mem[96] = 144'h07000981020f0ab600640a140d850cf3f02e;
mem[97] = 144'hfe4b00dcf800046d00d0fc15f56c0384f071;
mem[98] = 144'h0cbdf57f0f35f98df404ff00fb21fcd5f540;
mem[99] = 144'h0f5dffb70ad30d9a01fef3720a9301080703;
mem[100] = 144'hfecbf108ffd8fe71f095fe3602bd072ef856;
mem[101] = 144'h0c0c013e092404f3034af3e4f41afa25f4b1;
mem[102] = 144'hf93ef8a5f9def054f8d8033d096804c3f765;
mem[103] = 144'hfa5c08680f5e027cff81fb79f74a077df65f;
mem[104] = 144'hfd0ef857f2c80d1606680105067e076e09af;
mem[105] = 144'hfd0a06d30b16f3c60060f9cff1bdf48ff630;
mem[106] = 144'hf68af18405d10de40253fcccf1f504a90518;
mem[107] = 144'h0487fe9c020ef265f55e03590068effcfa82;
mem[108] = 144'hf079fe65091a050e0664fb08f72ffe4df644;
mem[109] = 144'hf66d06abf473fa7af53cf03ff7b10c2c0ba3;
mem[110] = 144'h00a209affe1afd640f46f4710455f75ff15b;
mem[111] = 144'hf5c7f674f321f00c0870f76d0f62f1d8f472;
mem[112] = 144'hf869f43c03b0fea003840e20f3bdf2450b2d;
mem[113] = 144'h017f0b3a0c0f0d400de607fd0e2109e60630;
mem[114] = 144'hf1b8efecf91b0122f2f70315f19e03030573;
mem[115] = 144'hfdf9fce7fd38082ffcb7098bf23600810adb;
mem[116] = 144'hffdf0801f84bf67508e6fcb20f3707eb08bd;
mem[117] = 144'heffffc8d07e00847f788055af0fd0aa40dd0;
mem[118] = 144'h0a0c0c8d050a07d30b78fb530bbdf441f99c;
mem[119] = 144'h019b0172f90efb4009e70bf50a7af7660a62;
mem[120] = 144'h0617065208ecfbb10f330128067bf39b0dfc;
mem[121] = 144'h07840b840760fbb109edf02e0c4bfbc9f5b0;
mem[122] = 144'hfb2bfa2fff3f07380df7fd15f4c1fbeaf483;
mem[123] = 144'hfa2ef975045ffbbeff710f49f4a005f202a7;
mem[124] = 144'hf400069e0466f0effd0a035df363f8c50a05;
mem[125] = 144'hf42f061c0cad0605fd94f1df0e1009ebf2f8;
mem[126] = 144'hf579096d0cd0f0caf967f5a2014105a9fc69;
mem[127] = 144'hf45df2bc06e4fb1507de0afff5def8e10195;
mem[128] = 144'hfe7d09150bfe0ed7fdb7f0c2fc81071cfd3a;
mem[129] = 144'hff1cfbd1f762f9f7fce801dd093ef29cfe8f;
mem[130] = 144'hf3ea04d502f4faac04ea07000a1c0d3f0cd5;
mem[131] = 144'h0ab90c0cfcdefaa3f1ba0c02f8f6f81e01b8;
mem[132] = 144'hf0b0084403e5fc04fb80f4dcfb26f672fcdc;
mem[133] = 144'hfdab08130fee0d330292f5cffcaa0a170dc2;
mem[134] = 144'hf26b0594001bf913fc83fc940730f7e3f723;
mem[135] = 144'hf5d0f214f280fe9bfe36f502f38508d801e5;
mem[136] = 144'hf8ed0e5202e501140da2fd4c02920d7cf7fc;
mem[137] = 144'h0cb0ff4f03c60a63f818f5d9f8ae0407f5df;
mem[138] = 144'hf6bef09f076c0a290df303000daa07c203c5;
mem[139] = 144'h04e3fc75ffd5076500f8f68af154fd21f281;
mem[140] = 144'h04ef001cf2edf46ff5c60179f2980d62032f;
mem[141] = 144'h06faf0e60cc6f2d3f713f435f8a5fc4901da;
mem[142] = 144'hfebb025c0e0bf315f11df49cff99076800ed;
mem[143] = 144'h04fa02bc070bf682fae2f61002d109ddf196;
mem[144] = 144'h0aa70c24095e0ba009f6092f093608f0f669;
mem[145] = 144'hf9520e0bff2d025501fbf9eefe35086f0954;
mem[146] = 144'h042efbd40248f794fc15fd0ff362f964fb43;
mem[147] = 144'h014006a90e7c0c2df45904b901c20b4a0af4;
mem[148] = 144'hf62702acfea007c80b270bd8f85afa5c0c5d;
mem[149] = 144'hfad80a9f08a7ff49fbb7f5ad0f16f994f343;
mem[150] = 144'h0d13fff00c0d0db00735fcb0f40905f3f526;
mem[151] = 144'hf6e00265fb7ffca001680a150fe505ae0d7a;
mem[152] = 144'hf461fa68fa30039df30101cafc53f27e0ae9;
mem[153] = 144'hffe0ff9d0ffd0e90f5a20d28ff2208b80917;
mem[154] = 144'hf6d6f381fc00f47cf4f4fd8bfab9f58f014b;
mem[155] = 144'h0445f9a0f2d70b340ab606930c08078f07bb;
mem[156] = 144'h0bdd051bf6b90fdf05c7f44802200ecd020a;
mem[157] = 144'hf911f25503f30c40049c050aff9b0abaf102;
mem[158] = 144'hfc1d013c0206fa8dfa60f814fe77f2650a12;
mem[159] = 144'h076efab4f3520ad1fdb8097f015d08d8f421;
mem[160] = 144'h00a5f2dd08160dbc0fe7049f0cf707a00115;
mem[161] = 144'h0295f077f958fb5df5ff07b3f581f772fe23;
mem[162] = 144'hfbd2fbf803a20159f372031ff011014cf30d;
mem[163] = 144'hf0cc0a61fab600cffc71f1b603be0a53f17a;
mem[164] = 144'h0cbdfbd7f82c0cd5fddbff8a02e0031bfe78;
mem[165] = 144'h091f01c50bf80bbbf87609c00c6609d70bdc;
mem[166] = 144'h0fc7fe83f236effef8ecfd62f2d5fbf90c78;
mem[167] = 144'h020cf62bfa52f486fee5f93b0817f50007f6;
mem[168] = 144'hf05dfd1103defd8df443059ef157f2b3f04f;
mem[169] = 144'h026c00890bb70ab3f9a10ca606e8ff390083;
mem[170] = 144'hfa88f6daffaa0645f4ed0cdbfa9509a60da7;
mem[171] = 144'hf578f0b500a8f9330ceafd16041bfaf20a77;
mem[172] = 144'h0e510cdf00b7f3e8ff2704030b640967fd49;
mem[173] = 144'h061a02d00c67fee4f318f5d400610b2d06cf;
mem[174] = 144'h0246091403610549fb8af594037409f50f69;
mem[175] = 144'h01040525f582f7fff939015cf106fdffff3a;
mem[176] = 144'h0ac8f246f1bbf8b8ff19fc90f58e068ff578;
mem[177] = 144'h024102af0799f3fc02edff15ff17f1f6f8cc;
mem[178] = 144'hfa0dfde501ecf35d03f5fd9ff89108c8094c;
mem[179] = 144'hf01df040f447f887fe9e0dfcfceff05a083e;
mem[180] = 144'hfc6effbd01190b8403610b8207b00f0effe7;
mem[181] = 144'h088201defaf2f2860f82f1cc02f6f091fcb2;
mem[182] = 144'hfd2f01640ec5ff11fc6b0a5cf2c401b808d0;
mem[183] = 144'h0cd900590409f508f3f3f1a8005bf7c109ab;
mem[184] = 144'hf0fa05890cc8f41ef1d0005c025e0939f43c;
mem[185] = 144'h0790fb45f1c9f2a8f3370ae30159f16f085c;
mem[186] = 144'hf8c40d6a06f10652f7aaf042ff26f04eefce;
mem[187] = 144'h06e6f2f3f8800517eff807c0048afcfb0bdb;
mem[188] = 144'h0e77fecd0323ffee0be3f2daf3d10a34f971;
mem[189] = 144'hf624f88c069f071d07980ebdf951f707f96d;
mem[190] = 144'hf331000a0c540c920291f678fc2200e10842;
mem[191] = 144'hfe66f394f80606ca00000e21f0c7fcb30e5a;
mem[192] = 144'h0618fe4a0fa20deaf98af144f3730fba03ea;
mem[193] = 144'h0db10113058e0f450a0903080d0bf29608c8;
mem[194] = 144'h096d0076f8e8f46103e4f3e60e19fa6bfee5;
mem[195] = 144'h0922f30d0640f55dfa98f1d9f83cff230598;
mem[196] = 144'hf34300def2ee0f25fc15074df29bfe72fbef;
mem[197] = 144'h050602f809b80560049b02a6fca00aa9f44d;
mem[198] = 144'hf862fa6ef424f45df8ef0738f627f6330bfb;
mem[199] = 144'h064e0e4ffd13f097f7fff607ff280f0b038d;
mem[200] = 144'hfb3bf01df82904cf039e0213f8d1f3940aea;
mem[201] = 144'h0ad2f64cf5a70389fb1df840f6660c0dfd5f;
mem[202] = 144'h077105e70f77fbca0985059d063902e2f288;
mem[203] = 144'h05d3025d0e4c0e92f6c805670549034e0da1;
mem[204] = 144'h017008a8f05002a0f933046d072ef750f3df;
mem[205] = 144'h0357f3830efc05b6f38cf2acff0d03d80ed3;
mem[206] = 144'hfacd0f33001d0c28f56bf827f08ef644fe75;
mem[207] = 144'h038af7010834f551063403f8089ef7cd01d7;
mem[208] = 144'hf646005af6bafe0ff107fd7bf0ea064bf9c2;
mem[209] = 144'h094cf649f9d8fc0cfda5040bfc7df918f32e;
mem[210] = 144'hf9a5f991f4d4f2da0d10fb300588f2f805f1;
mem[211] = 144'hfe4f014f0d7af15f0b66f7e3fd480e2b0bed;
mem[212] = 144'hfb27fe5301f5f4d807130157fbf8ffdffc35;
mem[213] = 144'hfc7e02160ef70785fc520654f090ff8a0931;
mem[214] = 144'hf846f5e402fdf90601ef0ce7fe0308e3098d;
mem[215] = 144'h0c52f3b80274fec1fe170597f89a0891059b;
mem[216] = 144'h09b5fdd9fc60087c0a62f2f2f9ceeff8f9ef;
mem[217] = 144'h04b2fa3d07fef6480147f6adffbbfbee09b0;
mem[218] = 144'h0694fbab0a74020d00270de7fb2af98b04a0;
mem[219] = 144'hf5b7fd09f21c02b8f833f58df22ff6ddf943;
mem[220] = 144'hf397f607f9dcf3aa0308ffd8f600025c01ec;
mem[221] = 144'h042ff56cfbf6f0ecf33ef775f04c0f550ac4;
mem[222] = 144'hf64604b1f6ce0be1f1dafedffea5f505f782;
mem[223] = 144'h057e0317f44ff823f44d09a3f6fdf53fffcc;
mem[224] = 144'hf17a0bd1087df4ae079ffb59fa28078c0c97;
mem[225] = 144'hf2f2f196fa85f13cf6ccfefffb86f6e70857;
mem[226] = 144'h0370ff4e0774f9f20365017efc57fe2205db;
mem[227] = 144'hf93d0b66ff99f576036dfc00fc39feadfa97;
mem[228] = 144'hf5b6f48e0b45f3f0fa1e042ff2c80f17fea8;
mem[229] = 144'hf79dff49f796fc51f3b50cee08b6f349f440;
mem[230] = 144'hfae2f3affc1d0138fc10090bfa3103dbf2ab;
mem[231] = 144'h07c80efeff4700fcf60805900ed20b210f94;
mem[232] = 144'hfdf00366f64b00c60305ff0b0077f08a019e;
mem[233] = 144'hfe5a091cf03102d4f2d8fb240541fdbe0df9;
mem[234] = 144'hf92d0fc80fe2fbe30f3a0457f7edf521feab;
mem[235] = 144'hf31af763f626f03a04a7ff76fe120583f3be;
mem[236] = 144'h098ef999f8f5f0c3fd78fc40f57200a307fe;
mem[237] = 144'h00a704170971f0350d0af39dfe41fcc4f299;
mem[238] = 144'hf79b045606790396f408068df5c8fb5b0ade;
mem[239] = 144'hfe0ffb60f38bf160043c0f36f8a8008ffbfd;
mem[240] = 144'h0aaff91a0f7efd68f1190f8f0b81f35afbc5;
mem[241] = 144'h0884f4baf3e1f4f60e81fe5ff54df4bbfbef;
mem[242] = 144'hfec8f033f1450a01ff87f4110b6cf0e1fd79;
mem[243] = 144'h0b9ff875002e0d9ff64efd3bf3150b320096;
mem[244] = 144'hf7f804e30747f6330e61f89cfa2e086a06f8;
mem[245] = 144'hf3ecfae2fd5704dbf9a3f91a063a025cff64;
mem[246] = 144'h09380295fc8bfa9ef40ffa760489f722f521;
mem[247] = 144'hfe3a0b79065b015c04a802a0fa34fba3f04e;
mem[248] = 144'hf49d0c6e0a1503b4fb80f560fafb0205098e;
mem[249] = 144'hf95ff1f607f30d990476fdcef3bdf69bff7d;
mem[250] = 144'hf034f20e0f1c03bdf2f2025c0b55f075faff;
mem[251] = 144'hf5f1fc1c093cf9c00e7c0b6ffb410cfff7cb;
mem[252] = 144'h08b6f89709670e3c08f50139f5360a18fe18;
mem[253] = 144'hf9d6f87ffb6df9cb00860f33f44f0559027e;
mem[254] = 144'hf8880ba109c0ff220608f81306b40d9b0529;
mem[255] = 144'hff06fe3500c60dd905a4f3f7f855f5540bcd;
mem[256] = 144'hf30707d2f4ed0d72f520f97efab504bc0b1a;
mem[257] = 144'h0524f0590a07fb8ffe2307fa0256026b06cf;
mem[258] = 144'hf957f575099e00620273f29b0571058604f2;
mem[259] = 144'h04fe08ccf01ef372f48af53af4210121fe6e;
mem[260] = 144'h047f0596013df83e0b3102f0fe7f0f5a075b;
mem[261] = 144'hf6a809cf0fadf06df1200b56f122f4a2080b;
mem[262] = 144'h0432fb72090c09d5f4b4f65f077ff2a0f09f;
mem[263] = 144'hf3b7f1a80d64f132f75df43efe490571f72b;
mem[264] = 144'hf9f202b3f1b6fa130f050712090a0e80f06a;
mem[265] = 144'hf2df033906b4fcea0074031ef70e069afb7e;
mem[266] = 144'hf9d5005d03630627fa66003c0c240a2cffa1;
mem[267] = 144'h0c380464f2e1fd2709c1fee4f8460eee084d;
mem[268] = 144'h089dff18036904040186f9610962063c0c81;
mem[269] = 144'hfadff5c609be0e1c01e6f8be0f3908a6fbd4;
mem[270] = 144'hff22f22c0556f10afd64f9e8f984ff1cf5c3;
mem[271] = 144'h0e790ff309b4f34bfba80dd9f554f47705f4;
mem[272] = 144'hff360eeef4ddfd37f078fa3cff0f0d460199;
mem[273] = 144'h0d510312fe2e0d72f57107b6fae1f5af0c98;
mem[274] = 144'h0a7ff97afcc50b7e0f32f92f036bf3600426;
mem[275] = 144'hf9130433f5cb0a8408570df70366fda8f58f;
mem[276] = 144'h0f2e07f5057d074d08d10baef502f664fabb;
mem[277] = 144'h03c60951034c02bbfbe1fce807790d600e6a;
mem[278] = 144'h07b5f23200fb008b068604cdfa920f2efa18;
mem[279] = 144'h0de309b1f98409b8f43106160107fd97fa61;
mem[280] = 144'hf3e307d0fe4602bef8330f63087ef3c7f9d1;
mem[281] = 144'h07040824f9ba0dc8f019fbfdfdd600e3fd33;
mem[282] = 144'hfab2098df7c2fb9a0f9ffc0c0ba006d0f784;
mem[283] = 144'hf883f4dffa9cfb120356fd25f16a0fbd001d;
mem[284] = 144'h06400f73ffa8049bf05cf471feaa026df983;
mem[285] = 144'hf1d8fc4b08f90ddaff060bddfd59021df66e;
mem[286] = 144'h0f33f6c400bef4450713fb1bf0b10f7affa6;
mem[287] = 144'h03aaf4e602f30d8503c0f44df004fe58fa92;
mem[288] = 144'hf5290b33f9bd019cf9c401850e2605e105b5;
mem[289] = 144'hf844018a0b1cf94d0261f2e3f1afefd3fb8a;
mem[290] = 144'h024007bf0a7d0f58009705a8fe01f64700c6;
mem[291] = 144'h04a0072508f2f4db04d8f40e04f6f0c00b18;
mem[292] = 144'h0d76f9ca0b8af725f9950d9ef1eaf103fedb;
mem[293] = 144'h02f3f8eef068fa8a07140fde09ef07250df8;
mem[294] = 144'h0ce1fa71fe66f5edf891f37b0a150490f683;
mem[295] = 144'h0313f8a3010704d4f1a1f09b08fd04c4f7ce;
mem[296] = 144'h0addfd0cf7cb0bdf0f1d0d67f849f2dafdea;
mem[297] = 144'h0c6408a70f1d07ac06f80ee3061908c4fc4a;
mem[298] = 144'hfe3407580e8bfc07ffc60bc7f5920884f997;
mem[299] = 144'h0dd4f6fa04080eecfa85054e0c25f40c062e;
mem[300] = 144'h08c1f1d3fd05064efa9b04f40bb9ff25031c;
mem[301] = 144'h056a07fff0b50478079f08c7fca3fec9febd;
mem[302] = 144'hf02a0e120d1d0af204740403f3fbfde70419;
mem[303] = 144'h06480f92f78209a60027f03f0853fd40f698;
mem[304] = 144'hfa5d064cf4a1f4700597fa0bf10cf538f8e9;
mem[305] = 144'hfe700302fdfc054504bcff85f0a1efff044a;
mem[306] = 144'hf23d02920f12fa67fb28fea00e8a00cdf611;
mem[307] = 144'hf86e0ca0038b0b63faf308090ade0023f17c;
mem[308] = 144'hf1b809bd01a9031a0bed0e6ffe38f509fc15;
mem[309] = 144'h0ee8f6b90e97f3aa08cb039af1d8f472fa17;
mem[310] = 144'h0fee02e2f0650c100aa40c59f7e9071e00e1;
mem[311] = 144'hfa84f07d059202d308abf393fcf80594fee3;
mem[312] = 144'hfe400baffbdd0d570187fd00fb7104c0f027;
mem[313] = 144'h048bf7990316f21d0633fa64fe77f4910524;
mem[314] = 144'hf65e031c0e86fb2ffec903a1f7060f16f278;
mem[315] = 144'hf988f96ff5b80b1afd120361fac30f78f8be;
mem[316] = 144'hf01cf34e0140faac0815f096f986fbc9f5a3;
mem[317] = 144'h062c0dabf73801b6fe49f282023c0b21f94e;
mem[318] = 144'h080405b5f99cf0a003bdf1c1ffebf035f156;
mem[319] = 144'h07b7015000a5074905dcf6b90f81f990090d;
mem[320] = 144'hf31ef73c09b508bef9d807200400093bfd35;
mem[321] = 144'h0fd5f727fb2cf8ebfa930d500373fffb029b;
mem[322] = 144'hf87b0647fd51f6d20f50fff60a4603e40028;
mem[323] = 144'hf593087b092a02edf1a6046fffe50bd00087;
mem[324] = 144'h0cd8f98f0d21f592fbfdf216f90e06fdf1e9;
mem[325] = 144'h0067f7d0f18d051ff30e0e95ff8cf68c0d50;
mem[326] = 144'h0f0affdff9f9f1acf544029303700370f0da;
mem[327] = 144'hf946fb2c09e306ec06850e680d030e18f54f;
mem[328] = 144'hf31704aef4cef932fe0707d4f89df6bdfe38;
mem[329] = 144'h00d00638fe40f463024b027c0dc2f8560ed6;
mem[330] = 144'hfba2f36304f20860fe650647fdcef9ae0c9d;
mem[331] = 144'h093b05ba0670f9e002800faff6850929f1e7;
mem[332] = 144'h09c0f9faf36b07a80576038ef8490bd1f13d;
mem[333] = 144'hfc690dab0ecc05000b3a0040f280fb2d02a0;
mem[334] = 144'h0cf3fa6ef98df67ff449081c0e46fa7601e4;
mem[335] = 144'hfe25f08500d1fb21fdac0c6e0072001f0cb0;
mem[336] = 144'h0fa4f14b005a0e0b0433f94b09ed088601c6;
mem[337] = 144'hf6ef0a27f226f37705f602b60faef8d70564;
mem[338] = 144'hf57709b1f1af00950fbef1dff051fbe607e2;
mem[339] = 144'hfbcbf69b0acdf649fd6ff9cff9d30cfdf76c;
mem[340] = 144'hf614f8c501d00268098c0e46f65f08dd0f72;
mem[341] = 144'h0e1bf6bf0ed9013c0d60f13d0fc0ffab03eb;
mem[342] = 144'hff2c08e4f89d012a05a908fb0b5c0f2cf4ea;
mem[343] = 144'h001e042406a6fcaf03c5f82df3d4001a0e26;
mem[344] = 144'h0e24029202b902cf0cc0fe0bffaaf7c201ac;
mem[345] = 144'hf605fa7c09c90bba09dcf4cc08ba007307e5;
mem[346] = 144'h07ea017dfcfef36d0f7a0e8ff172f8b00206;
mem[347] = 144'hf74c0a0fff25fbb4fb45fbcbf2a003290dca;
mem[348] = 144'hf1960828006804bdfe81f445f716f5d2f081;
mem[349] = 144'h006bfeae052e0d31fba30322f852fdfaff59;
mem[350] = 144'hf255fd9c008804e0fb3300f5084bf8b1f3ff;
mem[351] = 144'hfe4e0a44f84b0b5a00e1065c0232f03b0ed8;
mem[352] = 144'h0c9bfab1fb4d0959f7c5f2c00042fb190a8e;
mem[353] = 144'hff48f944f5550b6afdd503bbf545009f068a;
mem[354] = 144'h01ed0b43092ffb480cadf25af46e0367fd6f;
mem[355] = 144'h0133f16205fe0985febff3b2f56df9200ce7;
mem[356] = 144'h0fc3f8a70b77feaf0a23ffe4005004a30314;
mem[357] = 144'hf76201a1fd3cf5ab05e8f5a0fc6cf92a0493;
mem[358] = 144'hff480a48fcda042af7c00317f5b0f8040352;
mem[359] = 144'h0afefb8508c8f6cd01550e810bc5fe22fb93;
mem[360] = 144'h0eccf13101c9fd3d000a0b26fe70f5b4f7cd;
mem[361] = 144'hf82c0daafdbffa51f136046ff052fc7d02ec;
mem[362] = 144'hfa350c6cf3020559fad5f74c040a0c2ff428;
mem[363] = 144'h0a80f97b09abf625fcbb0b52fe1eff89f4f0;
mem[364] = 144'h0e1904e4f48a0e17f1980f320e07fde7f8da;
mem[365] = 144'hff8efa35f74df21bf1b60068f064fe980cd5;
mem[366] = 144'h0521025efc27f52e0cf2076a035bfdb6f129;
mem[367] = 144'hf71df1a9091c01dcfc2b080df2c5f9590b5c;
mem[368] = 144'hfbf60d11f8abff3efeff0a260efcfb71f249;
mem[369] = 144'hf923f22604ebf83b0162009e05650deffd31;
mem[370] = 144'hf677f3c404290b7f07bbfacfff730b150799;
mem[371] = 144'h0da5f4e9f29a093101220e92f18ff43f014c;
mem[372] = 144'hfa72086efe7d0c410ff7f22df09ffad1fe67;
mem[373] = 144'h01e400d20b3bfcaaf3a1f36106740534038f;
mem[374] = 144'hf2320cb5f75b0c260499f5950023f8fb0288;
mem[375] = 144'h0e42006b0b7c0406f0e2003d04d8f315f2be;
mem[376] = 144'hf8cd0410f499022d0d41fe400d490cd5029e;
mem[377] = 144'h0197003cf6fe0869fa41038b0da5f4300f4c;
mem[378] = 144'h0f4ef82af3580d0605bf0734f2f1fd3dfff2;
mem[379] = 144'h0f1ff528f34e0311f0110962fd06063805bc;
mem[380] = 144'hf4f2fd0dfcbcf08a0981f3330b43fd95fbda;
mem[381] = 144'hf0d0f38af414fcc00de10d6105e700bdf866;
mem[382] = 144'hfd2afeabfd630a07f250fee1064b0638fdf5;
mem[383] = 144'h062a08d206630af4f1a5f6e6fa01f138f703;
mem[384] = 144'hf0f006d802fe022b03f4075f0bc8fc7c0eea;
mem[385] = 144'h04cef8750e48f55903f5fc650b24f96e071c;
mem[386] = 144'hffc005080048f83f0545fac1028e066e05f6;
mem[387] = 144'h07f806fb09cbf30f0a7d0a2ff739f001f328;
mem[388] = 144'hf748fa31f523f035f171f4ea0a8f04f20f1a;
mem[389] = 144'hf2b0f9bb0c5bffba081df5bef6dff343f19b;
mem[390] = 144'hf9bf022905da07fcfa93f29306c4018f014e;
mem[391] = 144'h0b1e0fdaf8c00a0c0218fe07fdcafe4d0f07;
mem[392] = 144'h0b04fcb50f5208510dac06e60943fdce040e;
mem[393] = 144'hfa76f7defb5d0c2dfd45fae0f34af37701a6;
mem[394] = 144'h0eb6fca80ec20982fbc8f650026dff3eff85;
mem[395] = 144'hf7870a79046bff58058af5bf0fa9f1d50127;
mem[396] = 144'h0746f418fa1efced09830b4202370a810cb2;
mem[397] = 144'hfa23f19c0774f545001cf0d20664033205ea;
mem[398] = 144'hf032f0fb069a091bf8d40fbc0ea206ba0309;
mem[399] = 144'h0a9cfa1ffe610ae00fd10a3105ba03eb0514;
mem[400] = 144'hfa8c0efd030d0c3a066ff9b5f7a30a52f629;
mem[401] = 144'h0d3c0c9d0e32008afefef1abfee4f3c50b98;
mem[402] = 144'h0748080e02220ae207660f7ff927fc740e65;
mem[403] = 144'hf4b3f412f442f5740fe6f4c6fba3fa200b65;
mem[404] = 144'h0e28fb64f792fbbef78df96ef65ff1720609;
mem[405] = 144'h0a440a7eff4efdd907c10c0dffbf085a0542;
mem[406] = 144'h0d59f124fb8afbd3fec30a84f7260e5b0e8a;
mem[407] = 144'h013b06eaf5c202130eadf7e3f42809eaf814;
mem[408] = 144'h0c09f6c6077a02e1f39a050503fbfe5bfbbb;
mem[409] = 144'hf52df34002daffef0b4ff0cafcedf3a8081d;
mem[410] = 144'h0b13f8010d87f68b0914fe1804da071dfd77;
mem[411] = 144'h0e83fee2f1dbf58b0d5cfb69f47005320e92;
mem[412] = 144'hf4d60b84f9120db0078f050bf0e704d2f530;
mem[413] = 144'hfb530c0504b203820dbbf3bdf9dd09850e44;
mem[414] = 144'h035df433fef3fc070ecf0de00df4f1330b7d;
mem[415] = 144'h024805a9021efbc103f20c8b00d4f246f562;
mem[416] = 144'hfcb4f080f5b403a40d140df6fac802b20eac;
mem[417] = 144'h0a5efae30297f8170292f951f5880884ffd5;
mem[418] = 144'h0e8f0677f9e402a6fdf3080dfe0b024cf9da;
mem[419] = 144'hf017f710023c034afc3cfc92022b00f6f15e;
mem[420] = 144'h09f2059d0393f535fdc9f566fda60bc2ff9d;
mem[421] = 144'hf59df28bf2e304540a2a03aff1c7f96d0ee9;
mem[422] = 144'h05f50ea3f62a0b19069bf4e909daf80f0430;
mem[423] = 144'h00aa0bfffb2d068b0a8d0bc2f096fd36f191;
mem[424] = 144'h0400fed2f36cfd1d079cf227ff77f60af307;
mem[425] = 144'h0d2d08da0432ff1004940763f2280e4cf8a0;
mem[426] = 144'h02d7fd7e0b32020af1adfad9009df4d4fcb7;
mem[427] = 144'hf5e008690981f1740fc4f3330ae30fc0fc73;
mem[428] = 144'hf207f2f0fac10d7808fcf4830092fb8505a2;
mem[429] = 144'h0dda0169fae50ce5fb29f4b404b9f0dcf9df;
mem[430] = 144'hf6f400310e0af27700f0004cf917f48200a7;
mem[431] = 144'h0cb1f296f53c05fbfb1bf028f4e7f4ef0044;
mem[432] = 144'h0bdefa930a4108a1fbce0385f17cf4a70f18;
mem[433] = 144'h0fecf4adfc22056df347037dfe930329f15d;
mem[434] = 144'h085c033607ca0700fcc204b0fcb1f7cffad4;
mem[435] = 144'hf40efe720259fa56f605feca02300a68f475;
mem[436] = 144'h0d8df110fde1f2700b1c077f076bf329fb6f;
mem[437] = 144'h01fcfca2ff7bf4a7030f0830f114f4f70d56;
mem[438] = 144'hf90c0c8ef3a4ffbdfb5ef1e10268010d0311;
mem[439] = 144'h00c5fd710d6a0707fc83fc75fba602fff2e1;
mem[440] = 144'hfebb05caf2bf0d1f052603a2f9990d970784;
mem[441] = 144'h0ac40cb4f74d05e8fc9dfbb7072efa3e0afa;
mem[442] = 144'hf3770563f04d030df377055bf226fd23fe1a;
mem[443] = 144'h079f0c29fafcfc42f75c0dfbfa3afa470ad7;
mem[444] = 144'hfc3207040e920793f2860b280f3cfcbc08ec;
mem[445] = 144'hf8ab0304f63e05e4056904d30245fcb9f9bf;
mem[446] = 144'hf5f2ffca081706d803a7003cf6e607410fd6;
mem[447] = 144'hfade0067fd4c0c9d0977f3d3fed2f41df90a;
mem[448] = 144'h00310021f8e4f394f481052f0225f26e0855;
mem[449] = 144'h06ba041c0061f4cdfe550efefb78ff8a05c8;
mem[450] = 144'hf28ff135fa8dfaf2f6ea0c40f4640721fc29;
mem[451] = 144'h0d57fee1f07af8890fb9079808eb057bf6e1;
mem[452] = 144'h06fdf4cc036d0cd6fc5d0c2600db0e4dfdcc;
mem[453] = 144'h0a080cc103d80d8001f2014cffa8f827fd1b;
mem[454] = 144'hfdc4f4b0049ef41ff9bd02c60f360270f14c;
mem[455] = 144'h0400fecdfbee044d09e0f2e7f08cf293fde6;
mem[456] = 144'h062af89c00a4f5040877f78d0cc509550639;
mem[457] = 144'h058900aef095f94ffc1efdda0e3af1280347;
mem[458] = 144'hf6300d88ff4b011407b30f5c0c03f77207e1;
mem[459] = 144'hf6a6031c068af0740bd0f2340049f281f2de;
mem[460] = 144'hfe7af2480162f5df0a2407b90568fa76f4d7;
mem[461] = 144'hf9090e7b0121fe2df04503b80c9ef9f7055a;
mem[462] = 144'hf103fc75ff87fde3fc5008ebfebaf2cef1cd;
mem[463] = 144'hff0c039efe970b8bfff3fb7ff6fcfcfb06be;
mem[464] = 144'hfa38ffa6fa6cf5c6f9ea0a2602b6f364fe2b;
mem[465] = 144'hf701044a088bfee8f805f84ffe09fc050386;
mem[466] = 144'h0e03f6360c34f0250c3100610e66fad5f0c5;
mem[467] = 144'h0581f2cd0de6094105b00bec02d40d2f08d4;
mem[468] = 144'h0c22fd7df792fdb1f3ee0b3ef89cfc23f699;
mem[469] = 144'h0e5e0bef033f0ba80a2ef61df9660ef0fa17;
mem[470] = 144'hfbb20533f9cdfe930794fedd0c48ff42f720;
mem[471] = 144'hf8dff42e003101430cfcfa95fef2f3930389;
mem[472] = 144'hfa09061dfa27f499f4170105052af591fb70;
mem[473] = 144'hfebafe32057804f50586f3f40578fcb2ffd5;
mem[474] = 144'hffcdf5b001e8faa2fa28054dfa8af566fe23;
mem[475] = 144'h054d09b1f59005d7064afb79fa120762f9b9;
mem[476] = 144'hf327f8b10c0c0ef50158fa110b26fe3605be;
mem[477] = 144'hfb60fb9f0175fa240589f2fff0bb02d60dfc;
mem[478] = 144'h03720f0df1c40dfbf3b4f7ebf70809ea04b7;
mem[479] = 144'hf635ff730fd50739fa3b0c88fd8801d10cde;
mem[480] = 144'h06960221f351f9580e66f354f0ff0ea70c83;
mem[481] = 144'hf7430cc5f15df5a3f4ccfd2cfec8f8cdf561;
mem[482] = 144'h0f23fa63fa71f5ed0debfbf6fb83f281041c;
mem[483] = 144'hf39f0030037803b60dbf0f21f3860819fb35;
mem[484] = 144'h0ba7f6c80ddc017c0d49057c0883f41d0133;
mem[485] = 144'h04c4f7230257f8340e9c0825f211f690f431;
mem[486] = 144'hfffef1d1f22df3960907feb40870ff64fb40;
mem[487] = 144'h00acf2d4fd07f3d709b608baf4340fb5f4d7;
mem[488] = 144'h007b0e13ff20031e0f22f5cf06edf6e50858;
mem[489] = 144'hf1b5063201f80cc5f22b0d30fec40f53fdd4;
mem[490] = 144'hf2c20c820687f488ff65f4430e700ddcf004;
mem[491] = 144'h00a30a790d0b0359f2ae09dff03df93cf87a;
mem[492] = 144'hf8b40ecdfb4d06a2fb71f3aef55101f7fae4;
mem[493] = 144'hf684f302fa2dfb190ce00196fde6fa04f3a3;
mem[494] = 144'h062ef4530ece015d037e0d4206fa060407fd;
mem[495] = 144'h056807b908c40ce40b0e060df975083f009a;
mem[496] = 144'hfe300e6cf7c609c20ec6f46f0ac6fa5807f8;
mem[497] = 144'h091dfbcb05320b16f9e7016cfbcdf857028b;
mem[498] = 144'h036d048e0963003b0e5d0c470ac8f9a50209;
mem[499] = 144'h0ebaf270056305ed045807260480f558f0c6;
mem[500] = 144'hfb7008520682f2c9f5d5098d0e89fa030ea3;
mem[501] = 144'hf65bf77f057e0024f165f55806670cf807ec;
mem[502] = 144'hf50a0bc604a2f91d01000d000c42f94a0759;
mem[503] = 144'hfa91ff68f909f077fa340a780b0904e7fe6a;
mem[504] = 144'hfb0bfe6ef33c0a2a05680f70f69409590693;
mem[505] = 144'hf17f0ea8f29f09b103d9fa4ef4f2f7e1f5ff;
mem[506] = 144'h0dc105f0f9f5f861f29dfeaa0d1c026af7f1;
mem[507] = 144'h098309bafbe7ffe5f173f272075ffee8f985;
mem[508] = 144'h07030b54fd9df9d80418f9cffc1c02280497;
mem[509] = 144'h0b2d098ff1ccf601f7f6f9dc0eedf9640c14;
mem[510] = 144'hf98aff8affb305e0fd9bf2c5fbfdf1160f2d;
mem[511] = 144'hf87b067ff95d0cdb084af625f3e1f13ff247;
mem[512] = 144'h0fe40e14f404fcdff1b2f2b7051401c2f531;
mem[513] = 144'h01960762fbf60b35f9d608adf3d9079e084c;
mem[514] = 144'h0e75f6b80986f0bbf365f7ddf116f961fb7d;
mem[515] = 144'hf3baf542fd79061d04a703e4f2310eb40a75;
mem[516] = 144'hf4530491059c02d602e0f32df3910c86f5c8;
mem[517] = 144'hf26b0d9efc33ff73f51b0b7af9ddf4e3f9fe;
mem[518] = 144'hfe1701f30b15fceff6a3f4e8fa37f5c700bc;
mem[519] = 144'hf8920d8706f2025404fef1c80e6704220162;
mem[520] = 144'h0194f8780f06fc340bf4061d0a26fff702e3;
mem[521] = 144'hf84b03c70e8b06f90343f095f23eefec0bac;
mem[522] = 144'h0bb806d904560542fcc6f0b00e62f9a5ff75;
mem[523] = 144'hfcce05640ca702660bddf90cf3f00ea6f6c3;
mem[524] = 144'hfb5b0d1d07d60932fb9dfc60f24c0d00066c;
mem[525] = 144'h0babf6ea0418f5bafbf4f7bf07bdfade0667;
mem[526] = 144'hfcc201eaffc0f617081f01c2fbb2fd43f2ff;
mem[527] = 144'hf84df5e2f57d051d05c4f8eb0462062bfe76;
mem[528] = 144'hf6d6f02e077500390ca5069b0d490b970abf;
mem[529] = 144'h0b40ff6ceff60f850ca6feaff4d50c8bfa46;
mem[530] = 144'hfa8af24af165017ef1c2f53dfd8df0bafd6f;
mem[531] = 144'hffbd07e906790dcbfc390aeffbadfb09fb92;
mem[532] = 144'h09c60adefc98fd0d09fe00b9f0c508f108a5;
mem[533] = 144'hfbb704b2f117f1340a8b0a97090cff12f0ed;
mem[534] = 144'h0d41f9e2f33af23cfc4209620720f76b06a9;
mem[535] = 144'hfbe4fe270751fcecf37cf9c7f6420bb00b45;
mem[536] = 144'h06ca090f0868ff9df1b8f94905effa1cfa21;
mem[537] = 144'hf4e2f1380a1105fd05a80d9bfe980544f2c5;
mem[538] = 144'h060dfc4cfd460131f57bfba7f7aff3e803f0;
mem[539] = 144'h0eb60150f83905db0e7f06c0f3f2f0090125;
mem[540] = 144'hfc490f6cfcd5f9d8f27ef56a0de705a6ff7a;
mem[541] = 144'h01c6f17105f3f68afabb0bff009205aa0da1;
mem[542] = 144'hf05802e4028705e1f0e5f8e2f4f00950f96d;
mem[543] = 144'hfd9fffd1f5800bd6fc970bb2066c077d0420;
mem[544] = 144'hfb7c013e008d0e6ff7480b0d0dfcfd99f517;
mem[545] = 144'hfb4e0e2f070c0b26f9b2fb2d0d200d13f237;
mem[546] = 144'h0cd60f5bfce1f8d2f53d0513f24af57dfea8;
mem[547] = 144'hfb8ffab3ff0cf3d6f0e1fc17f92c031d0931;
mem[548] = 144'h05cbf6a604b8039af85bf1e0fd81f62d0acb;
mem[549] = 144'h0f7bf8d4f2a9fccaf01b07c8f5910dc40720;
mem[550] = 144'hf2a9f31ffacafc48030e056cfe9aff6affad;
mem[551] = 144'h0f8af9d8fefa0d3b0a640a480765f8a0f77e;
mem[552] = 144'hfb89fd5e0c4ef838ffa20573071ef22801d5;
mem[553] = 144'h04ab08f0f1d003320f3c04d1fccbf88c0844;
mem[554] = 144'hfa3e0a5e0430fa0dfa39fa92f6930621f8b6;
mem[555] = 144'hfe5dff4df710f0c60ea403450d91008d0445;
mem[556] = 144'hf2d404b6010e0914f16a08100f09f791023f;
mem[557] = 144'h0adb0946f53bfc58f1b6f6acfdbc041afd0b;
mem[558] = 144'h0074fc84fa150f7a0fa604e7f517fa000a0a;
mem[559] = 144'hfaa3f22903320def0289fa39f60bf98ffc7a;
mem[560] = 144'h0e32f617f303eff904d6f9c9f08902a3f2a8;
mem[561] = 144'hfe390c79fdf1f13706780a3ef708fec700f2;
mem[562] = 144'hf002f69d0ee2064700e1f82efa0a0b8cfa0f;
mem[563] = 144'hff0af9c3fd15036b02fa0cc207b907670c26;
mem[564] = 144'hfdcdfe06fe60f14a0f8b0a09f20ff5900d10;
mem[565] = 144'hf8f7f3c40fb9fc1c050b0714f0c7f45805d9;
mem[566] = 144'hfbe8f1b3f6c5087a09e00d6807ad05430969;
mem[567] = 144'h081bf7d0fb8cf3b8024c00a5f1c7054ffb91;
mem[568] = 144'hf56a038e0580f6c4ff9d025e07e007b3f6e8;
mem[569] = 144'hf61c031d0eaf049f016dfddf0c9d021bf026;
mem[570] = 144'hf96903f0f7bc0b20fc630dab00170eb5fa88;
mem[571] = 144'h064cfa02fd86f6eff40b0f9800790cd50f00;
mem[572] = 144'h0ec5f904f5c80c940503f46e07930ec9f577;
mem[573] = 144'h016c06ab011c0ea0f4b3f2360d7ff437f3d1;
mem[574] = 144'h04a40b43fa1ff272f984fc2ffc6af29c0d9e;
mem[575] = 144'hf71ef8ae0ac5005e0bd8083d049a0d83073e;
mem[576] = 144'h03a9ff8d0257f05806a7f9fdf2d705b5058e;
mem[577] = 144'h07c8f5500c690140f4e00a3604ff0807f00a;
mem[578] = 144'hff770f76fd420c2df23bf50b0e1904d4f700;
mem[579] = 144'hf1e10a340fa2ffa507660933f2230bdd05a4;
mem[580] = 144'h0e4e076d0fadf188fe1efb0ff4040c96042e;
mem[581] = 144'hf744068ef858f53f0b15009508a308e6003c;
mem[582] = 144'hf1790edbf2bd0db3f2d901de01bbf121f667;
mem[583] = 144'hfe400e150ae3017ef8b1078c003ff231fe3c;
mem[584] = 144'h04cdf5c00a4c027702790a2900cf0e81f4e1;
mem[585] = 144'h08efff000619fc18fa7107e7014c084af278;
mem[586] = 144'h03390a9c086dfc780877fa1100eef178f36d;
mem[587] = 144'hf1c1ff7b02fff451075f0748f4b70cdef4ce;
mem[588] = 144'h0424fe48faa8efd10dc10e680152028cfb0c;
mem[589] = 144'hff5502970f27f752f8bf0506f9f906d1f4c8;
mem[590] = 144'h0a7df012f71f0046f471fe05f70bf6d20796;
mem[591] = 144'h0fdd0fdf0978f5bdf9e2f669fe1b02e0031b;
mem[592] = 144'h053df0ab04b5f621fd0cf771f5cef0e804ea;
mem[593] = 144'hfe660afa01f204f3f27bf9be0c1a037a046f;
mem[594] = 144'hf4b5037bfa93f0bbf036f8d10b240b36f3b4;
mem[595] = 144'hfa8e0f5dff8700f104e60d080832faaa0172;
mem[596] = 144'h0e70f35af2fefea3f7350a86f2f308a402fe;
mem[597] = 144'hf453025ff1640b5efbe40d05fcfd050e09bd;
mem[598] = 144'h0a42f2e0f81b0dfc085af669fd000e4a0e27;
mem[599] = 144'h0b00fae1f536f7d9f2e7fd16f398f19b0c8a;
mem[600] = 144'hfac7f7ccf70a09e90d12f7eaf119f0c300f5;
mem[601] = 144'hf736f78ef75c03830467f1eaf834f561f416;
mem[602] = 144'hf869f2b3ff3df6fafdf6042ef16806910893;
mem[603] = 144'h0046fde3f5f7058a0f3606d30c49f1350db1;
mem[604] = 144'h098bf257fd62f3b00d89033e08880c94fe3a;
mem[605] = 144'h0461fd68fa09ffdbf4400888fa8b02190074;
mem[606] = 144'hfd71043bf4aaf2170ecdf14d0a8cf47c021d;
mem[607] = 144'h0a4f0eef0b7c063f03380ce6f35ef3930815;
mem[608] = 144'hff1c05530e200125f697feae0cbaf2d90216;
mem[609] = 144'hfebd0ab40c9506da04850c46faa403cdfb27;
mem[610] = 144'hfa02f7b60421fad3f2eef98ff588f893f424;
mem[611] = 144'hf8710eeff3bcf712f1dffd5cf7a2fe9b0c87;
mem[612] = 144'hf100fe39fefc0a39f5e90732f75d092708a4;
mem[613] = 144'h0ccaf3de075b048806d7f8c1ff5e075d0c87;
mem[614] = 144'h09a304c5f662f9c10bc2f7fbf1ddfe1d04c5;
mem[615] = 144'hffef0b92fbaff565f6f9f75f04890b8ef8b9;
mem[616] = 144'h00a40c2809a5fda207fdf770fed5f657f9a1;
mem[617] = 144'hfeacff470061f25c066df6f0ffcd0dfb0dc7;
mem[618] = 144'hf9cef0a8fabcf29205f40729f1390b9dfed5;
mem[619] = 144'h044501ebf216fd29fb9e052dfcb4ff100df4;
mem[620] = 144'h04d301560226f6b1fcec0cdc06dff71c02b6;
mem[621] = 144'h093b076af301f4c60cdafabffd000f64059b;
mem[622] = 144'h0183060b00e40572ffd900d00b010796f13b;
mem[623] = 144'hfc10f0980b7c08b60c49fad9076cfc4bf1c5;
mem[624] = 144'hfe0ff141f23e0ae40b16fc110b7f08370722;
mem[625] = 144'hf2b9fee3007b0397078cf195fe94033af810;
mem[626] = 144'hf57a00930b74fd7c0370f03001220c7c0e48;
mem[627] = 144'hf7de026e0b7507ecf4e3f22cf75ff548f32f;
mem[628] = 144'hf8d6ffb20632065c0657facbf6c2f6d5f8bc;
mem[629] = 144'hfdc8f543fb5c0099fc4ff358f7e4f5990f8d;
mem[630] = 144'h0af7fbbf038a048c0a5f03d5fffdfd8ff7b8;
mem[631] = 144'h01a60dbb03b80d98f443f47ff5240c3bfa4b;
mem[632] = 144'h03ecf456f84400100c52f8830622f511034b;
mem[633] = 144'hf85508160e6df6b2fc490828f755fdeb08a2;
mem[634] = 144'hf944f057f43df3e50fb6f69a086b07ba032c;
mem[635] = 144'hf984f8430511f3b8004802e8f926f43a0fc0;
mem[636] = 144'h0b5df6a3f4e8faf208fff201f9b1fd980e83;
mem[637] = 144'h09b408eaf7bafd68f3ddf9d7f03909cffb85;
mem[638] = 144'hf8be0cae0732fb010f1707110a74060d0985;
mem[639] = 144'hfecc01bd0a7cf3760e8a03c3f578ff5dff37;
mem[640] = 144'hfdbdf5c701bcf0190932f64b01c004a707eb;
mem[641] = 144'hf0360bd704930c02f96a07b40b38faf7f2c9;
mem[642] = 144'h02ed06a908fef270f1a4f74ef96af690ff94;
mem[643] = 144'h0e4ff75ffabef81a07fe0d07f05bfeb2f2b1;
mem[644] = 144'hf220062f0e2001990bfff6b80373f61bf01a;
mem[645] = 144'h01e306fb083b06bf0d8dfb3afbeafbc1fcd2;
mem[646] = 144'h050b01c10c4b0d3e0d41fbd1007607bef8b3;
mem[647] = 144'h07b1faa7f5f2f3c4f5dff8e3f1f40f4506b6;
mem[648] = 144'h05acf90207b4055ff58bf6d50986f67bff20;
mem[649] = 144'h0882fb0c0ef8f9cf0ca2f744f53af1880155;
mem[650] = 144'h0c9709b20416f878f32afc1dfedd0ee4017b;
mem[651] = 144'hffd5f367088905f3f9f3f70dfbf40428ff86;
mem[652] = 144'h0c3700c6f923f1a800bff1c5f8b60d9306da;
mem[653] = 144'hfd91f596fd470b250806fda9f6df0a0b0b62;
mem[654] = 144'h04e8045601a8041e0b0e0176085c08aefe72;
mem[655] = 144'hf09d0de6043cf0ab0c920e63f6620e770976;
mem[656] = 144'hf360fb3a0dbb0b7bf72506eff7c0f51bf22a;
mem[657] = 144'h05830aa0f2fd0895097cfe3b0c24014903d9;
mem[658] = 144'h0506f836012ef259050f05710cb80eb507cd;
mem[659] = 144'hf108f94bfa15f64dffca036df422fe8bf0e8;
mem[660] = 144'h0a6e0dc80435f66d089bfadffc9a04a8f896;
mem[661] = 144'hf064f0bd08eef26cfedcf38c0ab70674f762;
mem[662] = 144'h0e950b0006c50475fce3fb6c0058f7a1f2f5;
mem[663] = 144'hf89ef886fe850973f4b8f90001ab0c920238;
mem[664] = 144'h0d7ff75afc70081bf2230f18fe94f9d001ff;
mem[665] = 144'h0ab70cf708b20c20f2c60b29fa1afcc00961;
mem[666] = 144'h0d52f313fe870a6dff64f39a059c0de705e1;
mem[667] = 144'h0b950ec104730443f3dbf59cf9b50c38ffed;
mem[668] = 144'hf97b0b480cf709090e6dfbdaf572038507c5;
mem[669] = 144'h05dd00aff7d8f021f1ec0e5cf5d4fd52fb17;
mem[670] = 144'hf2780608f354fb8c0fb1f3a9099a0b5c0db9;
mem[671] = 144'hfa1904d50981fd38f951fd8f0796f54dfcd5;
mem[672] = 144'h013d0bfbf069f53bf88509680c030e58045a;
mem[673] = 144'hf5b1f92bfd910f21051c089e017bf41b046b;
mem[674] = 144'hfb2af3ab07bbf250026d0f69f29afd42f9f3;
mem[675] = 144'h0cff058ffc140be3fc4c0802f6b3f417fa5f;
mem[676] = 144'hfcaef4f603bf046af85dfeb20741f38f0115;
mem[677] = 144'hff47f883f0e70daf00c803630c2cfd38f462;
mem[678] = 144'h032109790baff5de0c45f0ea003307c405c5;
mem[679] = 144'hfc5c00d507d3fae0f8e4fd63f49ef41609c6;
mem[680] = 144'hf2c6f884f05b008ef89d0e35f29d0b86f485;
mem[681] = 144'hf9aa04e9f198f67ff136f5ba034f0b9e0210;
mem[682] = 144'h008bfab7f118052b09f7f4210317f583009e;
mem[683] = 144'hfd1af237042e08e80a2af17e092808920c47;
mem[684] = 144'h06f1feca0894f2990756fc1e057e0b84053f;
mem[685] = 144'hf9a6f56ef78af321f2740da0f6470d96f4b8;
mem[686] = 144'h06140b1f0c6ef33705080e580c22f91809d7;
mem[687] = 144'hf17d0885061c03b500dbf2c006e4ff0fff6c;
mem[688] = 144'h0be7f7c20886f2330d3900f104a7fb0df463;
mem[689] = 144'hfe26f1a0f0f1f699ff5306ae09fa088afa76;
mem[690] = 144'hf1b1016d076f0c93f251f831092df750f00a;
mem[691] = 144'hfbc702460b9ef0a5f8fe026cf6cd044bf514;
mem[692] = 144'h0289f1a20492f1730f8a00e50eaf0016f6f8;
mem[693] = 144'h0aa90eb0097df0c9f0d5fb46f7bdf7d5fdc6;
mem[694] = 144'h0bfa07070a990af7ff1c0856fd5bf8f00d8e;
mem[695] = 144'h08150300096ef3260544f100fbc3f4e801ee;
mem[696] = 144'h0058f068f4f7044df6910c7e05c60038fed3;
mem[697] = 144'hfcfa00d300a3f82ef84df94cff0ff1740ca2;
mem[698] = 144'hff9dfceb00260de3f20205a700e106aff47e;
mem[699] = 144'hff5d0fceff040cbe079c03a7079ef3910618;
mem[700] = 144'hfa1df5daf1d5f5520d4204f8f51ffb5defff;
mem[701] = 144'hefd0f00e094d0da0f8fbf3adf8d1f84b0d37;
mem[702] = 144'hfa79017bf5f2f6b4fe3707f5f41c029e0e30;
mem[703] = 144'h0a1bf2b00de80668f879f816f585f7870fb8;
mem[704] = 144'h0a190c8c0e170a5ef1b1f0b8f9b40f0606fe;
mem[705] = 144'h098bf1c106830f6c02d7075f066704b6f177;
mem[706] = 144'hf175f6d8fe110ee0f79e03cdf5860a000388;
mem[707] = 144'h052ff64b00e9f115f5d80fcf0cee0c840fd5;
mem[708] = 144'hfaf20371f4d90710f168fcc907f105cf0d33;
mem[709] = 144'hf1cdf0a10cfaf6f2f6e0025d06410c100aa0;
mem[710] = 144'hf1840210f0640f23f0eef77104ccf1bf0219;
mem[711] = 144'hffbb01dd05c8fb3bf353fda8f66309d00b33;
mem[712] = 144'h030bf332f53ff36cfa7cf1130a3e02b2fcc3;
mem[713] = 144'h0dd302a002570a7afa400fbd08c1f15e0ac5;
mem[714] = 144'h0c170f96efde0e2b03f806a50e7f02a1fbcd;
mem[715] = 144'h09800dde08b904d302ebffa3fea5f198f3b9;
mem[716] = 144'hf8eff2ab0f93082508df02dff9020176011c;
mem[717] = 144'hf0210dd60a48f91af6fffa9e070d0e040eda;
mem[718] = 144'hff5f0223097b0ef1f73ef98d0cabf9040919;
mem[719] = 144'hfa340994f05c0ee90ae1081bf642f574f811;
mem[720] = 144'hfec80bfa09b2f9620976f7f0fefaf1adf8ec;
mem[721] = 144'h077af5f00564f98a02d40abbfd630146075b;
mem[722] = 144'hf1c9f9fd0b36fc85fb3c0f1906e1fb5cfb71;
mem[723] = 144'h0e840ea8f0cefe040e50f541f8e3fdadfd4b;
mem[724] = 144'h0f14f7c6f7d4fd93fb03080ff285f506f39b;
mem[725] = 144'hfa4109740e9b002609e6039cf867060f05d2;
mem[726] = 144'hf0bbfc39fa9efa580e6f054d06fc03920d27;
mem[727] = 144'h0547f3f2fb470ba9ffb0f1a5efd3008cff1d;
mem[728] = 144'h07a90496fef0f6bc0515f98a0e010260fe58;
mem[729] = 144'hf6710303079efe1c078ffccd0a46f9df0aad;
mem[730] = 144'h03b80f6af088fdde0c53fcdcfceefbb8f68a;
mem[731] = 144'hf1a20171f1dafc8d026f034b099cf94b0758;
mem[732] = 144'hf7b9fd30043bf5e6023602b6fe160182f4f3;
mem[733] = 144'h0de9f4e403220f3cfc8cfddaf9f30ea2f515;
mem[734] = 144'h051c036202180463f710f871fc64ff8f0b9e;
mem[735] = 144'h01ddfc37f4d80686032b09a60b1b034e0b9f;
mem[736] = 144'h007b06920b9af7d60ab509aefa91f5230a34;
mem[737] = 144'h050f0cb00ae80fdd04a00abdf24809bd0ff6;
mem[738] = 144'hf2440f11ffbafa08f40effbff757fff30493;
mem[739] = 144'hf303fabef7f1f214fcb306aef30df5920808;
mem[740] = 144'h034f01dd019a0081058af0dc0bc6fbf2f885;
mem[741] = 144'hfc4f08dd0dbef451f3510703fe0a059af987;
mem[742] = 144'hf6630bd7f190f7fd01a507e0052cfbf40450;
mem[743] = 144'h0cc501eb00dffb5af2020e0009d1092b08ca;
mem[744] = 144'hf58b0614fbf1ff62ff5cfaf8f37cfeb205f8;
mem[745] = 144'h089804800a870e600cab0e0bf8edfde8f621;
mem[746] = 144'hf4a3f6f502d4004e0a9ef03309b2ffedf0c5;
mem[747] = 144'h00790b35f0f1fbf9f8280c9700840ada0a03;
mem[748] = 144'h0a7ef6f40f5af46df404fbe302c507b8ff88;
mem[749] = 144'hf3ae0f17f4abfec500ff0667f687f93c0f61;
mem[750] = 144'h00360565f7a6f8a40dd4f53ff730f1620f25;
mem[751] = 144'h0097f1b100fefce90b30ffaf0c7003e70509;
mem[752] = 144'hfe99f4c9f03cfd13fb1c08c0fb88f0950757;
mem[753] = 144'h0e2802710bf7023a0068f13cf391f37a0251;
mem[754] = 144'hf080f9e40e5701b407a9f9a2f6a007ec0b12;
mem[755] = 144'h05eef4ca07280f57f473f555090cf96f062f;
mem[756] = 144'h055d05b6f7b80d29f1d0fbfdfb9b09deff5a;
mem[757] = 144'h0741f31c0c57f810fe1901d4f314f0fdfbe4;
mem[758] = 144'h027c07e305850232f917074fffcb0a330f1a;
mem[759] = 144'hfab2ff21f9a00dd301180e320ce503760fcf;
mem[760] = 144'h01af0fbcf6ae041df6c5f6da0dd5f23df7da;
mem[761] = 144'h0423f42204dc02e307c00fa0050afd6404b2;
mem[762] = 144'hf38efbd706c0f1d5fb43fb1c0fef0aa2f735;
mem[763] = 144'h03cd0343f123f6fcf20f0be4f1fb060105ab;
mem[764] = 144'h00fc0d2a0e3808400125015bf335036cf0cc;
mem[765] = 144'hf824fff7004e0d74ffb9f213f6380ed1f354;
mem[766] = 144'hf877fad3fab5f85f02a00bbbffc503f1fd69;
mem[767] = 144'h0edf09600e500ea8fc50fa5df82c06cf0db7;
mem[768] = 144'hf6380faafcc3029bf49d0ca4084105ef0498;
mem[769] = 144'hf4a00c050426fc700a300acffceaf42c02e1;
mem[770] = 144'h0f280e4709870958fe43031bf6ea0a9ef33e;
mem[771] = 144'hfd32fa82fdd6041f0152f289055cf1e108a9;
mem[772] = 144'h0ba0feed002107fcf1bff5f909810d190526;
mem[773] = 144'h0ef306dc0ac10d0905a2fe62f99204b1f5ae;
mem[774] = 144'h08aef229f79e0774fcc50a0ef313f19f0465;
mem[775] = 144'hf975f8a10f47081701940249fe19088c0189;
mem[776] = 144'h06290bb3f4650bc50a980f7e075bf65af771;
mem[777] = 144'hf7eff902fcb5016f00d1f948f3e7fe8ff25a;
mem[778] = 144'hf4b8f624f7750bd8f53d025d0406f70cf7da;
mem[779] = 144'h040afdcdf413fbc3fdfa0d980c1e0dfcf804;
mem[780] = 144'hfd83f1c6f46bf5bb000dfecf07aa0026f4c6;
mem[781] = 144'h0bde0e23f5bb0c34f87ff14503ee0cd704e9;
mem[782] = 144'h00eff6d0065400330590f29100910d15f08d;
mem[783] = 144'hff21f4b0f821f8df048cfff70c4f0ea5fc34;
mem[784] = 144'h0b8af25a05410d55f276f9fdf12000940d60;
mem[785] = 144'h0640fe38fb58ffc4f094f220f0ac091a0ad2;
mem[786] = 144'h0783fd23f441098bf09001630f40fc9f02d3;
mem[787] = 144'hf393f39ef85d0500f0f9044a039bf1ec0d31;
mem[788] = 144'hfd71051109a30ec90213fbe7092af5240ac0;
mem[789] = 144'h0f0cf17c0d240130feb4faf20ed9f1c9fb58;
mem[790] = 144'h0be8f151ff2d041efa2d07ae09eb0c2e09a0;
mem[791] = 144'h03c70f7cfe2a049b0ab908a8fbb40e19fe95;
mem[792] = 144'hf0c0f13a060bf580f711f9ccf9bffcc6f40c;
mem[793] = 144'hfc680b39fc0d057c0ec00cd1083bf61d0cab;
mem[794] = 144'h0edaf5b9089efa4c01470108f8020e9ef5b0;
mem[795] = 144'h0113f1db0199fba201aefcd8f85df9600b7c;
mem[796] = 144'hfd3b001e070c0e02f6400b09f425f3770d6d;
mem[797] = 144'hfd3d08fb003dfd740e0ff293fb86f6880104;
mem[798] = 144'h043afb080a5d023106870d3df7f80755f67d;
mem[799] = 144'hf2a3068e03ba076ffdf0fcf6f83e038b020b;
mem[800] = 144'hf08ef770f4210a030997f1d10cc709df0792;
mem[801] = 144'h08c1098c0383f5f10f230e71f92e0b7ffe37;
mem[802] = 144'h0810f029f7690b7505c9f427fc22f2dd026d;
mem[803] = 144'hffbb089af601fa61017901a4fafaf0aff9cf;
mem[804] = 144'hf25109dc053b083c04d4fa8ffa920794044e;
mem[805] = 144'h040bf1df01f20b3df071f1d8fd410765f7f4;
mem[806] = 144'hf2670b06f188f0b408ea046efc6ef25d0be9;
mem[807] = 144'hf5d1f699f8db0cdffe99f94ffb8305040b55;
mem[808] = 144'h068d063a04fd064707200682012101b70168;
mem[809] = 144'hf832f606f1adfaaef7eb0aa9f0b3f13e0615;
mem[810] = 144'hffa903a2f788ff940804f7360be604470a37;
mem[811] = 144'h0ca3f9eb0700fbfc049cf315f7cbf013f99a;
mem[812] = 144'h0a3707b20efcf66ff6bdfa1208c2ffdffe5e;
mem[813] = 144'h0842054b0763082bfd71f58d06e40826f012;
mem[814] = 144'h06f8f281f89906f905050216056207f10ce5;
mem[815] = 144'hf91a0e46ff000d0bf485019bfdfdf71b0ce6;
mem[816] = 144'hfaf10f7b0e4c01120fbdfc24f6510f5205ae;
mem[817] = 144'hf2fdf9ec0de4f5d3fff9fc500567f47c0572;
mem[818] = 144'hf110f9ecf41609880c2f01ab0454f87e00b2;
mem[819] = 144'hfec5095cf6ddff37fcb008b60617019df68d;
mem[820] = 144'h0be20b67f12dfe04f795f0970e6601c809d1;
mem[821] = 144'h0b4009410c3100be0618fe350d820f81fc4a;
mem[822] = 144'h0b3302c80ae5f977f02ef32bfbe80ac20e9e;
mem[823] = 144'hf6c9f7ff05a5fab204f4f2fcf936078f0790;
mem[824] = 144'hfc14f332f73c019f052bfe790609fdc90187;
mem[825] = 144'h0cb1fa22fcd30f7a0214054dfec7041cf670;
mem[826] = 144'h042a0e2f05600344f8ea0f5df1ce026f0343;
mem[827] = 144'hfc28f023f39307fefdd506baf00b06cd0b85;
mem[828] = 144'h0716fbeaf33cf91f03c901840a960343ff67;
mem[829] = 144'hf8c9fa0dfa4ffd89fc4e0945fcf7fda60c2d;
mem[830] = 144'hf5fcf400fef1f7f50f790a3af1be0d3df6a3;
mem[831] = 144'hf56e030a08ad0a44020df6770cd4f8abf505;
mem[832] = 144'hf874035b0946f2c9f75905400f4008cbfdc8;
mem[833] = 144'hf4adf0cc00eb0baef2ec066201c204f0f71e;
mem[834] = 144'hf3c3f4f70117f034f479f4c5f17d0956fe8c;
mem[835] = 144'h0c1002c9ffd6f0850859f1c1f7790204f255;
mem[836] = 144'h063a06bff6a8fe93040f05ed0a82f6020251;
mem[837] = 144'hf93d08cdf6a70b0bf732f6fe040c067af641;
mem[838] = 144'h0dc605240327f3da077b0ffbfa130646f9e5;
mem[839] = 144'h09cd0e6dfefbfcb20f2e0be20ab9f805fba3;
mem[840] = 144'h0ea909e0fb170dd1f7390e1cfc32fee0f30f;
mem[841] = 144'hfcbb08d7f69ffd02032404f9f7f30976040e;
mem[842] = 144'hfca2f518f49802f70a0bf7adf65ffe350698;
mem[843] = 144'hfbc308160cb9fc47fd520dda064ff9890fc9;
mem[844] = 144'h03240234fce90f3708600e500f300b3ef3db;
mem[845] = 144'hf50bfb420a95f6500791f28d0dc8f933f3f9;
mem[846] = 144'hf2d60bb2f2200ec1f8b909a7fdf5fa150398;
mem[847] = 144'h02f8013208f7002c072f035b010ffe37f90f;
mem[848] = 144'hf4b5f95efd2609ed06baf7adf275075d086e;
mem[849] = 144'hfb8bf341f86b04c0fa71fbe1fb7b0098f9c1;
mem[850] = 144'hf8590fc6f1c60d5809f2f846f75f0df50ee1;
mem[851] = 144'h0520f288f10cf666f533f179f9d8f9ba02b6;
mem[852] = 144'h0aecf86dfce6005e00f6058304210614ffbc;
mem[853] = 144'hfc0d0f7108f7f774f6c30706066807a3fe25;
mem[854] = 144'h011602adf8ddf472034cfd60fcf1032a0341;
mem[855] = 144'hf36d07b507f70623070efb310f1af2f80dee;
mem[856] = 144'h0352f22907a202c207a5fc2107c80d42fa29;
mem[857] = 144'h0bde00fb09b80e9a05d3f7dd071701d1f079;
mem[858] = 144'h09520b0700c3f99507c9fee60da9030400db;
mem[859] = 144'hf3a60e700f2bf49df186f599fd3efd3dfd61;
mem[860] = 144'hf9fff9e1f6e2ff03f37c0dc8f892eff6f7b1;
mem[861] = 144'hf917fa9f04ca0c59fb55fbb40f60eff3fa7a;
mem[862] = 144'h09c00a4dfaa0f5a9f2fc09180ac809190b76;
mem[863] = 144'hf4550a8d00c2f954f758f142086bf1830152;
mem[864] = 144'h0e67f2fafbfe0a1006970e0af6e7f15efc1f;
mem[865] = 144'hff07f9fafed10fe00754fbfaf056f01deff8;
mem[866] = 144'h0c96fe68fefef093f81700eb0bfe022ff5d5;
mem[867] = 144'hf8e5f62cfbec0b78fefa02a3fb6f0824015c;
mem[868] = 144'h05a3f9790d62f77900750aa8f975f99809a5;
mem[869] = 144'hf75e0e3efd6cf3cdf29707c501be0289f2b4;
mem[870] = 144'hf1aff83e0ee10773054ef26e007d0070f8c6;
mem[871] = 144'h05ac005ff947f7d004b1052ff6db08cd05bf;
mem[872] = 144'hfd7204aff3410e140c8d0c7a0e2efeb8f576;
mem[873] = 144'hf363fb7af5b1096a033ff3920b3d069609df;
mem[874] = 144'h060f07b3f6b806edfea80446fe74f9dafc18;
mem[875] = 144'h0e590f040790f2bff51d02cb0a39fa370f13;
mem[876] = 144'hf529f95f0390f89f062604b70fcf09350e23;
mem[877] = 144'hf801fd0a05b0fb5bfbcef933f43000cbf9ed;
mem[878] = 144'hf92ff21e089405e6036a0f4dfba4fbe2f705;
mem[879] = 144'hfb6e0c4cf400fb92f16a020ff432f4f00052;
mem[880] = 144'hfa32f05dfa16008bfab9fdedf47f0ee7f602;
mem[881] = 144'h0b42f4d40a0ef80609680103069f0648f852;
mem[882] = 144'h0f0a01590f59f0ddf0c70a07fe8a0dd701b6;
mem[883] = 144'h050608cbfb69f22902e3085cf6de05690479;
mem[884] = 144'h0671f5f20374fe110673fdf603b70438fe1d;
mem[885] = 144'h0f65073b03f7047c0116f848fc090e26f829;
mem[886] = 144'h0c2a058cf29afe960abc07a5f8dbf7caf23f;
mem[887] = 144'hf60afe570812f9e6f163fb7f051f0669f1c6;
mem[888] = 144'hfb81049f09e90beb0715f7d10bbef6c60b1a;
mem[889] = 144'h05270cf5fc320e59f9b10e80f1d8f714f04e;
mem[890] = 144'h06bafc33000708bbffe40fd008d70b9fff88;
mem[891] = 144'h0d800a2ff34206ca08da0e75f4af00f90be9;
mem[892] = 144'hf27ff1f6f132f12df1e4f1950eef05ff0894;
mem[893] = 144'hf33ff5290f2b0ce70198f8f8fde80baff403;
mem[894] = 144'h02b80214fc1d07caf75a096c07b70113f1ad;
mem[895] = 144'h0087fb9ef94c0ae1f8040e370de6f24004de;
mem[896] = 144'h0ae102d3f826f77c0b020245fc4b02b9fd6e;
mem[897] = 144'h0786fcd2007f0fc8056d0f9e0a0e08410197;
mem[898] = 144'h0fc2f84905b706a000f906fdf00702fc03e5;
mem[899] = 144'h04a3fb43f8c9f9eff2abf5de05a00e000301;
mem[900] = 144'h0ca5032ef6fcf49dfbf504570f96f779f18f;
mem[901] = 144'hf0310e730f9af33102c6efeffe75f2dbfef2;
mem[902] = 144'hf4f20c6cf14700e3f2a70ff3ff0f066cf498;
mem[903] = 144'hfbcef9aa063806680303f547fe0b06500d2e;
mem[904] = 144'hf125064cfc42fbacfd01f3130fd2f87ffb25;
mem[905] = 144'hff80f209f86efffefa5809900541f2230ad8;
mem[906] = 144'hf3b5f83dffe30f76f5010ac6f846fa7cfa65;
mem[907] = 144'hfe6cf289051c0083f487043df1fd0013fd69;
mem[908] = 144'hf4e8fad9f22a07ed070cf459074608aaffa9;
mem[909] = 144'hf9c3f595f0f6ff710e0df8500709f6de0d4e;
mem[910] = 144'hf22efcfa048df5500c340060f167ffe80224;
mem[911] = 144'h0ee6f2c0fde4f78ff176fe2800130d690164;
mem[912] = 144'h050cf1d90309034ef008ff0d06c30f0406dc;
mem[913] = 144'hf93509b6fe66090cfd60f8ccf178fff40827;
mem[914] = 144'hfb150c250ba300fe0dba0000fedc0f66f0ba;
mem[915] = 144'h0cb40ab9f8420a57ffae00ef0788ff6efe2b;
mem[916] = 144'h02ba08d6fb2700bf03a60541faf3ff990f69;
mem[917] = 144'h062ef421f456f8a5f1d808de0d050d36fd8d;
mem[918] = 144'h0941fbfb037ef8ff06020160f0c8014bfa2a;
mem[919] = 144'h014306a9029400a8ff7e0380fd31f70ff593;
mem[920] = 144'hf593ff08f970fdf306a7f6bff756f02000a8;
mem[921] = 144'hf36d08b0f09ef37ef4f6f84505a1fcbbf4e9;
mem[922] = 144'h0dbd090300c5ff470ebbffc00f8df9e5043b;
mem[923] = 144'hf7b1fb710a4f07d60cd40be3021d074d0d9e;
mem[924] = 144'h08b10f5e0d3cf793f7cc0f44055df848faa5;
mem[925] = 144'hfc42fb85fa52f08604da0d89fd86fc88f9fd;
mem[926] = 144'h0145037af9350ce6f43bf5d8f199fc1708a1;
mem[927] = 144'hf73ff18cf04302bb0593086707def47d0b31;
mem[928] = 144'hfab30f2df2e7f85401560be0f108f5fc0eeb;
mem[929] = 144'h06c4fd0ef5b30118f1900b03fb880ce3f225;
mem[930] = 144'hf92cf314ffa700c0089c0c9a0a4c085a0470;
mem[931] = 144'h0c2bf44107d1038c08b40256f0390067f506;
mem[932] = 144'hfa64f30ff892fcebf9d5fb5ef77b080907f7;
mem[933] = 144'hfbfb0524fb84f2e4f5c00f8b05b5ff9ff0a1;
mem[934] = 144'hf9b4f9e00ed80adcfaf202f0f4680c310193;
mem[935] = 144'hf7d80cd4f90d0f3ff5ccf2980b120d4cfebc;
mem[936] = 144'hfcb0f3870b1ef7250e15feccf4b20a38faa3;
mem[937] = 144'h0523f7df02a501ed031a0004f0f3f9dd068e;
mem[938] = 144'hfa4dfa2609e100f7f2f1f64f0312081b0d89;
mem[939] = 144'h002cf830086c012902ddf0b6fb2ef91ef1c0;
mem[940] = 144'hf0e2f42e04c80cf0f102faed07d8fe8a0a09;
mem[941] = 144'h0696ff3ff456fba20444065ef3ff03b40869;
mem[942] = 144'h0c94091afd7bf7b60cb8f6cefd9c0b290857;
mem[943] = 144'h0623fec4fa7f08300b98fdb0f6e0fb7bf1bd;
mem[944] = 144'hf10f06710884f734f2980b4f04c40da1f767;
mem[945] = 144'h01a401bff648fc250bf6f158f021f4b1f52e;
mem[946] = 144'hf5f60a47f930fff9fcf20e6c0bbbf5b50aac;
mem[947] = 144'hfab60642f42a0d1af430032efb44090f086b;
mem[948] = 144'h0fc7fd14fc53f1c0f2f9fa29eff603d80284;
mem[949] = 144'h06c8fbfff052f8eafcf3033cf399fa69f4ab;
mem[950] = 144'h04a8f4d1f3cff4d707dcf4bff392f412f577;
mem[951] = 144'h06edfe09f297fb760c5f0e53ffe1feb8fb5b;
mem[952] = 144'hf79f094c0213ff9f0db209e0fc3a0d810c55;
mem[953] = 144'hf2320b86f76f047b0279f1acfe8cf7f0fbba;
mem[954] = 144'h0f1cfc1408df05b40d1df10dfd4bf813043e;
mem[955] = 144'h0c12f4cb0db004230c23f26f07cf04bc06cf;
mem[956] = 144'h0b4504350398fe960389fc3104730a4df516;
mem[957] = 144'hf84b03bcfac904e90553f904076df1a1f1c9;
mem[958] = 144'hfd21f628032401a2f08ef6f70a85f818f9de;
mem[959] = 144'hfcaef0f6fcfc03dcf11a029df5910c960fe2;
mem[960] = 144'h0026f92c03fff8a7f6bef8f0ff8d00fa09a9;
mem[961] = 144'h01bb05bcfefa0c87fdcdffe50c5ff6e0f410;
mem[962] = 144'h07c1fd9ff5d2f20f06f4fecbf997007afc95;
mem[963] = 144'hfda6f61309ae0c460660f14bf7a502400f6f;
mem[964] = 144'hf6a404330c1afba8053606120d16f7edfab1;
mem[965] = 144'hf40d012500580d08f53ffb77fbcc0b5f0507;
mem[966] = 144'h0bed0561fbcef0b2f431045d004c0bb101b9;
mem[967] = 144'hfa3a08b3f71203bff4e20403f74601f4ff3c;
mem[968] = 144'hf40109ebfb1e0a56021c0481f263ffcff39b;
mem[969] = 144'h06fefac3052104ea0a22fd3ef3daf423021d;
mem[970] = 144'h00770e640337f291f376026e0de1f41603d4;
mem[971] = 144'hfd43057c0e7608fef1a607a80cef019dfbf4;
mem[972] = 144'hf4f6ff93050f06f7009406130e76fdf2f640;
mem[973] = 144'h0f210bbef132fc36ff03f3db0b59f5fcf3b7;
mem[974] = 144'hfcb9f9ad0d90f319006e0fdafdeef4dafa70;
mem[975] = 144'hfe5e0c9df86e0f1b0955f2bc06b4051b0442;
mem[976] = 144'h037900190b2c070f0d0bfe170ef30c8c043a;
mem[977] = 144'h0e850b77f22efcc2f2e50ac00accf03f0102;
mem[978] = 144'h06fa0d730ec2f75cff66f933f78d047bfdfe;
mem[979] = 144'h09b8fcb2f9bdf7d80a95f8a40dae0887f494;
mem[980] = 144'hf928087d01c2f327f0eaf0d7041404e702fc;
mem[981] = 144'hf27b0dfd03c400710c3a0ec30b1ff0d702b8;
mem[982] = 144'hf4a50102f8c1032b06f701790e0b0f63053f;
mem[983] = 144'hf134022d0bcb0c2afea5f8f206c90460f0be;
mem[984] = 144'hfdbb044600a8f53cf10a01de006a05100ad3;
mem[985] = 144'h01930d66f132098df6f1f8e4fe6301a10e90;
mem[986] = 144'h0064fe120dd0f3750882f763fbb7027e076d;
mem[987] = 144'h06e5f15ef6c3f401fee90a3cf2b9ff5cf421;
mem[988] = 144'hfb6402880e77f1e1f049ff3df4def1fafebe;
mem[989] = 144'hfee7f648f814f633000af80d0b6af564f5dc;
mem[990] = 144'h0869f7820f94f445ffc80cc80d9d002905d3;
mem[991] = 144'hff34ff56f220f6fe0ef9f55a0d6a040afd41;
mem[992] = 144'h054a095a0cb3f7230d1efb350de00866f1a4;
mem[993] = 144'hfb9c0af2f3def1650f2300e6f13c09ef0903;
mem[994] = 144'hf60100c307faf39bfe100da30a900baff27b;
mem[995] = 144'h0d81facbfad50e89003cf5ab08630d540a41;
mem[996] = 144'h0a99006ffa5e0384fc480e020915fa6f0ca1;
mem[997] = 144'h02210c75f47ef8270ce60bd3f8b1f6c6f5af;
mem[998] = 144'h0b9b09c8f3e80490f0aef8e6fb45fbcb0128;
mem[999] = 144'h09ebf341f63900e10e52fffafdc405e9f511;
mem[1000] = 144'h0f96fa37f9e00ceef1c405bef250f99ef893;
mem[1001] = 144'h0f7efbd6f5220a2ff582f8c00ccef9f003c3;
mem[1002] = 144'hf39dffad04bdfd64ff77fdae0291f41f0280;
mem[1003] = 144'hfde2f11805e002d4f35df8cdfe97f8aaf92f;
mem[1004] = 144'hefe20334f815f0220aeb00adf4d708450e7a;
mem[1005] = 144'hfc400aed0291001df9d3052a02e1fe610e24;
mem[1006] = 144'h09ee0b44087404f50bbb0b16f49709a5f80a;
mem[1007] = 144'h05e9fdbcf1f90f8f0b4d01a6f1990e950378;
mem[1008] = 144'hf2c30b3f04c1fc39f17ff2c6f974f3290b39;
mem[1009] = 144'hf32dfc8df0b6f10bf7bc0cb7089f0dabf0ac;
mem[1010] = 144'hfde20bdb0e650f910e26ffe1fdfb031b0281;
mem[1011] = 144'h0bbc0d860519fe79f02600cefc22f6b70c22;
mem[1012] = 144'h08a5f17f04c0f726f24e040c07f5f3d00af9;
mem[1013] = 144'h0ca5f721f339fabbfd8dfdb3fdfeff4bfaf2;
mem[1014] = 144'h0b820044fc21ff6cfccc050c0dfdf5ff0be9;
mem[1015] = 144'hf173fcd8f0def3c502cc0660fd35f21708b2;
mem[1016] = 144'h01850008ff880b25f5e5fa720d04f47bf794;
mem[1017] = 144'hf1e80d730105f5a8053c0d93f088f9b8f1cd;
mem[1018] = 144'h048df1e0f2d4f9e90e2cf26bf5b800d10c2b;
mem[1019] = 144'h04b7f2720d8105370ca1f51d08020780065b;
mem[1020] = 144'h0bbdf8fbfac4fc95fbbcf1ba0c890dd00e53;
mem[1021] = 144'hfbb3053403800b78f3d501090a7ff31bf5fc;
mem[1022] = 144'h01180d4401750f53fa730074ff7df0c309d9;
mem[1023] = 144'hf9c30825f6bdfc320ee3f39c07b702390fea;
mem[1024] = 144'hf57bf8d1fd76ff3bf8ff0cacf656fca5041e;
mem[1025] = 144'hf9ebf153f369fc390d93f92c0dc9f29c0c68;
mem[1026] = 144'hf16cfb3a057bf24102850c1300030fc70be4;
mem[1027] = 144'hfffc0ad1f13f0c6ffb6a077d05dd0370f241;
mem[1028] = 144'hf66bfe1903880294f957f45203bc05010bca;
mem[1029] = 144'h037bf2980e76ffc0f430f4bcf9fd0c8c03e2;
mem[1030] = 144'h07daf5d4f9f80fc30b440fcff99cff4cf299;
mem[1031] = 144'hf963fa8b0aa209ebf7fb09600d940f2800a8;
mem[1032] = 144'h0029f436fe38f2b7fc05fe82ffe2f743fb0b;
mem[1033] = 144'hfef1fbd70386023cf9f8f8580d0f04e0f666;
mem[1034] = 144'hfaa8f9e4f2560b7afd720c39031d01210484;
mem[1035] = 144'hfb72f6f1f59d031a0e80f330f4390a1dfb4d;
mem[1036] = 144'hf027f64105090fddf88408a0f708f03e0bd1;
mem[1037] = 144'hf3e504350de5fe6efc0b08ddfb1c03f002e8;
mem[1038] = 144'h0929f93cfc44f3120c19f05ff1dbfd9e050e;
mem[1039] = 144'hfba400980dc40e97f87b082a09fbf91f0430;
mem[1040] = 144'h0fc90c5dfdbffdf6fb86016af6d5f282f952;
mem[1041] = 144'hffe9f6de05eb0f350810f771f46504b7f0a9;
mem[1042] = 144'h04f6fcc0f5b8f1af08eef6cef5edf41ff669;
mem[1043] = 144'h02b104220891fed90ef60d51065afee4ff13;
mem[1044] = 144'h087408faf2d3fa93f6d20e02f5d70e36f31a;
mem[1045] = 144'h09c7f6dc0cc00923fff104c5f40107220082;
mem[1046] = 144'h055708e60b52004b0a46004af730fe01f0b2;
mem[1047] = 144'hf9b6f844f3a9fdeb08880053f4b3f1f4065b;
mem[1048] = 144'hf999fccf09300dd001fc0549f49901b4f525;
mem[1049] = 144'hf163f6af0135f32a06cc07fdf9dbfceaf224;
mem[1050] = 144'h0f78f3df09290067f660fee801d6f881f85e;
mem[1051] = 144'hf44b05d9fd69fe8409c50f34f2e6f8aaf3b8;
mem[1052] = 144'h097bfdcdf2080dae0940f6160b75f194f993;
mem[1053] = 144'hfca7fd4f0273fbfafea8fb5606000e110ab1;
mem[1054] = 144'h0ff6fe04f23d078cf557f1d6033cf78003a0;
mem[1055] = 144'hff1d0c0ff35900bbf90a0cb0f71ef4cfff95;
mem[1056] = 144'h024c008efe7af0b20f550f140f5df442090e;
mem[1057] = 144'h0af500d5027cf64304910e41f171f3570159;
mem[1058] = 144'h08ca02e6f90f051806dff3a9f4a2f92cf2f3;
mem[1059] = 144'h0d820ba3061502b8f498f0f902c10388078d;
mem[1060] = 144'h03b50fb7fbbc07e3071afef80ace0aae092f;
mem[1061] = 144'hf0e6058d0964f7fe0974f52004430b9a0add;
mem[1062] = 144'h0d9d0cba0946fc40faacf68cf371f5190502;
mem[1063] = 144'h00f0fead07dafda40d31f2c4f07df8cc05e8;
mem[1064] = 144'h0200030301460e9f0563fa5d020b076b09bf;
mem[1065] = 144'h0eef033df21c09d2f46804270b00ff73f059;
mem[1066] = 144'h0f43f068fd56030c04ed014c02670286f377;
mem[1067] = 144'h00860b5c08cbfeeffa94f13809a80029f3a3;
mem[1068] = 144'hf8b0fd67fa6c071dffb602980bbdf2630a62;
mem[1069] = 144'h0ad70e80f8fd051d0e1df792f2e50be20297;
mem[1070] = 144'h0f12ffb50941fdfcf68af0110f7b099501c8;
mem[1071] = 144'hff5cf06dfe9008c0027cf5b105ce0f14f1fa;
mem[1072] = 144'h0f5707d1fd1f0e4908bf0747f09df15d0537;
mem[1073] = 144'h009e0a190058052b079504d5fb290423f5e5;
mem[1074] = 144'h0b9c0d2bf1dcfb02f48cf3fa0d04ff42f603;
mem[1075] = 144'hf550f6eb0dabf05f08ca0a5f0ec9f67f077a;
mem[1076] = 144'h0edb0b2d0e140902068f0ddc06e9f4affcfd;
mem[1077] = 144'h03cbfdd8f2d303cb031ffa360642fcfef337;
mem[1078] = 144'hfc93020803f4017104db043c03530d85f563;
mem[1079] = 144'hf3d8026c073df4a6fcdd057dfd91febb0931;
mem[1080] = 144'hf9fb0bd3fd440e490cf5fbcef318f576f22f;
mem[1081] = 144'hfde4f734f31bfa30fff4fabcf227f344013e;
mem[1082] = 144'h0e4ff450f78bf6860a21f3b5fb2bf7820d78;
mem[1083] = 144'hfc54f60c03c3f4d9f8ab0c3f0968f00105ce;
mem[1084] = 144'hf1370776fe260e1708b1f779f117fd15f85a;
mem[1085] = 144'h0e570087f006ff8df3fc0460fab8fd41fbf9;
mem[1086] = 144'hff78019bf06d0c4ef463ff1ff2ae081cfd1c;
mem[1087] = 144'h0f310ad0f82ff7e005fefe7ef46304d70aa6;
mem[1088] = 144'hf78a0193f9770d52fd13f31afc9c0232ff9c;
mem[1089] = 144'hff3c07af0df306c90d7607f4f0c3f953012e;
mem[1090] = 144'hfe72fb080dd5fb67f841050e03710f46032e;
mem[1091] = 144'hf69a01b9f758f37cf4b70683f520f0ee02cb;
mem[1092] = 144'h0d84f5c5032cfbda0fd1fca2072a09ef0952;
mem[1093] = 144'hf45806730bf10546f5ef0d7e03affb1a01f7;
mem[1094] = 144'h00f7f6aaf793fb130ec7f9f10567fa070091;
mem[1095] = 144'h02ccf93df48c04220c4efa4a0602007dffbb;
mem[1096] = 144'hfaae05b00643065a01500542098e036000a7;
mem[1097] = 144'h080ef6810aeb0d490d37fc480ac300100517;
mem[1098] = 144'h01a90f4afb8e012c0138f7d80c55fd03f942;
mem[1099] = 144'h04dd09fef178fdb40f180bb6f2b5f1170e4c;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule