`timescale 1ns/1ns

module wt_mem5 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'hfc0001d5ffe3face04250005029ef6f1f28f;
mem[1] = 144'h0967eb4aff7fecb30710007dfaa1eace032c;
mem[2] = 144'hf179fecaf89e0d52fce3ff21070ffca7ff1b;
mem[3] = 144'h084cef8c025f0a25f525f1f00663f7bf04ae;
mem[4] = 144'h0d74fa01f99af3c3f4020c3af1eafdc30bbb;
mem[5] = 144'h0231edd401de010ff645f930ee82fda50572;
mem[6] = 144'hffcf03400ce7fb6203aaf5db0319028f0552;
mem[7] = 144'hf73e02cfeebb03be0336f7cff932fa7cfacb;
mem[8] = 144'h0168f17f0603f6ec02430a0a03e4039c0d98;
mem[9] = 144'hf717fb950815f793022aff5df8ceede907c8;
mem[10] = 144'h00d0f992ef01f361f940f0d70a3a07b80364;
mem[11] = 144'hf0f4f1a7ffedfc5607740bd2f0a4f720fbb3;
mem[12] = 144'h01a2f376f9c5f345066d03d3fb2d0a58f829;
mem[13] = 144'hf46c02d8f9b9eeea045af978065202f6078f;
mem[14] = 144'hef41ff8b01e104710aaaf22207950ad9f4cf;
mem[15] = 144'h092ffcebf0fceffd04bcf705ee8df6c7f339;
mem[16] = 144'h003ffd86f8e5f8e8fcd3fbdc07b709e00cdb;
mem[17] = 144'heeddf31df360eb9507b303c4fe1e08fb0787;
mem[18] = 144'hf9100aec041efd14060efccb04fdef93fc9a;
mem[19] = 144'hfd4002760339f09ffa65f77ffe0d0725fa5a;
mem[20] = 144'hffe6f5d1fb2a039200e4f1ddf93a097dfc15;
mem[21] = 144'hfafffe30f8b908ee0496f42fecf1f25ff79f;
mem[22] = 144'hf4fb0cc0f3aaf4f2fbc0fb5cf930f742fa4a;
mem[23] = 144'hff3effc8f3a20b3bf6adfbaceeaa0744f98d;
mem[24] = 144'hfb31063ffeda048e0db30cf8ff930c7bf20f;
mem[25] = 144'hfb2af1b40996ee2001760a5cee59f60f0d2f;
mem[26] = 144'h01b90b140a210bb70079ef0d0999011e0a76;
mem[27] = 144'hf88404ddeeee0156f0dffa8a0830084604cd;
mem[28] = 144'h06270d36f7c8fb3a01b00344fcec0a6d01a3;
mem[29] = 144'hf1ca02c9f71ff836f0a40a4bf5acf786fca8;
mem[30] = 144'hff6ffbe6019a0481f0bf06f30cb4eff6037c;
mem[31] = 144'hfba6f61ffe1aec8406ca094e05d2f379ed09;
mem[32] = 144'h02be0db2f7dd0bc8f51cfb3aff3bf20bfbd7;
mem[33] = 144'h099204ee0bdeee46fae8fa4d0270f968fbb7;
mem[34] = 144'hf49807a4027d05e6fe8509d40500fb9c0309;
mem[35] = 144'hfd92fff7fa1f02d4f986ec7afedcf330ffc7;
mem[36] = 144'h086c01e5efc705edfc2dfe9cf68cf094f75b;
mem[37] = 144'h0014fec8084ff4ea07b8f46af1760814fd50;
mem[38] = 144'h069a04ce09c3fc91ffdc0248041302fa0982;
mem[39] = 144'hf331033afbccf321fd8dfcc10708077cf288;
mem[40] = 144'h011b0caa0d18f60d0ae8f458f88c0811ff33;
mem[41] = 144'h05b3f9d90576fad6f7f0fb7907700d57f18b;
mem[42] = 144'h0368fbdaf65c094c0b64075bf86504caf7fd;
mem[43] = 144'hf07eff1f07acf777002d071ff48cf537068c;
mem[44] = 144'hfc120517fbc509400d17f4a8fa69fee3f88d;
mem[45] = 144'h04a00199052ffa190b4900edf4d0038cfcbf;
mem[46] = 144'hf13e0746fd4700f5f6500a32005401e7044d;
mem[47] = 144'h08170494f80a057f0cf107aefd49fe64f642;
mem[48] = 144'hf2f50a160c2df43701ad0171f8b3009cef53;
mem[49] = 144'h0380f7990ae00c56ff89fbba0184ed71f768;
mem[50] = 144'hef11fad9f0760d8dfea10541047f06cf0479;
mem[51] = 144'hf6220dd7097c05d304700b3cf310f2220d1f;
mem[52] = 144'hf258f1bcf5dc0485f54e0492fb0ef6050679;
mem[53] = 144'h03adf1b50110f04bfc85028af7cc069200bd;
mem[54] = 144'hfca4f43d08c704a2f68c0a4f0c440300fb79;
mem[55] = 144'h03f60b8b0592edc7edab0c7d066b0691f380;
mem[56] = 144'h0790f9edff66f8a8fcd8faf5f70a06420b2f;
mem[57] = 144'hf1de09030d34facf0376f1af0a190d7102b5;
mem[58] = 144'h0d37069ff0dfffb7f020fcd1036e0193fe39;
mem[59] = 144'h091c0f3a0e2805ba0ebd00770de7f3d4f1a0;
mem[60] = 144'hfd3d0bb1f1abf7d703defeca01780d07f280;
mem[61] = 144'hfccbf283fe5a0918eda5f6faf86e07f8003b;
mem[62] = 144'hf6dffa8c02e1090cf703f89af083f2e10cc0;
mem[63] = 144'hfc4d0bb9f1b1f44802d70334eda4f00ff89a;
mem[64] = 144'h0aaf01b8fe3c05e402f8f847fb88f26000a2;
mem[65] = 144'hf289ee59f34d0117fd2bf3770344086b064f;
mem[66] = 144'hf40c061e02590fb1f41c0550fc69fd1b01b9;
mem[67] = 144'h0748fb860b0e08f505a30a0f08ec085b020e;
mem[68] = 144'hf3cf06e20f2404d605fcf9d203a0fdc9fa8b;
mem[69] = 144'h0fbc05a0f4a80db2f2e70eadffcff05df1b3;
mem[70] = 144'hf252fc7705db01a5fd5eff860633f09002e7;
mem[71] = 144'hf6f70db1f9bc0e2b0a15fb3608b10a880fa0;
mem[72] = 144'hfa4708d2062f0936f6db07740360f72306e0;
mem[73] = 144'h07fefb82f5cbf7c1f2db0cb305d70876f734;
mem[74] = 144'h08490ad309f5f620f8dbf0e6f95f03e2f12c;
mem[75] = 144'hfddcf1920e9702a7fb82f35ffccc00b70b16;
mem[76] = 144'hf8c6ff0b006dfbc1fdc6ffabf084fa38f94d;
mem[77] = 144'h01dff4eafd61085f0f600d900854fc6a068f;
mem[78] = 144'hfb46ff35f554091e0e30004c08c3f590f842;
mem[79] = 144'hff5e00a50196f6a8016bfc690c25f339fbf4;
mem[80] = 144'hfb91fb790841f7d1f4d00f60fa7200a3f7c6;
mem[81] = 144'hf06d0069f334fb030c3ffc68f4b7f3f0f891;
mem[82] = 144'h0463fc98feecfc7bf74c076ff7250d43fd5d;
mem[83] = 144'hfd4af902ff07013af08d011204210de5f234;
mem[84] = 144'hfdcafb8ff919039c0541f0d90db00e6706ed;
mem[85] = 144'hf061fed8f52808f2f0f1f4edf3260001f2ec;
mem[86] = 144'h0aa7fe25fe90035a051802c90ae00be6f182;
mem[87] = 144'hfc1905850e710762f5a0f6adf4770872fa31;
mem[88] = 144'hf6640c5bfc78fa1bfe250847065b00510774;
mem[89] = 144'h0dc3f51afdbffb13f7c00a44f6b60226f544;
mem[90] = 144'hf837f8ceff200185021cfb5e01a6f69a09d2;
mem[91] = 144'hf9090c70fb41087cf9a905a502c4f281f397;
mem[92] = 144'hfc9cf187f28df130f57af1b10c06f18f0f59;
mem[93] = 144'hf221f36b0c5ef8c7f65f0b93040d036df972;
mem[94] = 144'hffe60c7e08ad0ff9081ff33d06b40b1af065;
mem[95] = 144'h0d58faf0f49af45a0292074efb13ffbe063a;
mem[96] = 144'hfd39f42a0cd0f1e9f1bd06f5f72c0665fa76;
mem[97] = 144'hfe250eb8f01501e7fb1df2c000270ddff77b;
mem[98] = 144'h07d7f415fbf80a55f5b00427f42bff11f388;
mem[99] = 144'hf3c9012afbd9f303f74001b7f2380956f52f;
mem[100] = 144'hf4a6017c01380bf6005306860db3f2b4f0fa;
mem[101] = 144'hfe8106c3f818fa290044076ef84ff3f40e13;
mem[102] = 144'hf80f033cf27d0931fd55f9defbd60cfbefe1;
mem[103] = 144'h04140dc40151f9d5f0d20548f0d5f94ff57c;
mem[104] = 144'hfae204f1fdaff9140405f2020375f4a6fa18;
mem[105] = 144'h0f57fafd0f34fe44069ffde5f5fbf1c3fece;
mem[106] = 144'h05d0f147040c098afe6101fd0d3a08a805b6;
mem[107] = 144'h09490f78f89900fbfdf1fe3608eff75309df;
mem[108] = 144'hf77d016a0caaf7750218fc67089a08d9fe0f;
mem[109] = 144'h0dfa0a0600320434f436094e0c75f7150744;
mem[110] = 144'hf923f45df003041909b00e030c46fe0103c4;
mem[111] = 144'hfda0f9270d1507d60ce4f4f400c3f13ef52d;
mem[112] = 144'h004905b30154f8cffcc2f402fd2a0a63f092;
mem[113] = 144'hf95e025708600f430774fd04f52108bbf6d2;
mem[114] = 144'h09a3045f081f0e870581fedef5840d1c019a;
mem[115] = 144'h030efcd0f2650c580d2cfae004fffe750056;
mem[116] = 144'hf32ffb73f0660942fdd90ac20fedf086f7bc;
mem[117] = 144'h009df938ff66035f0022101dfeabf9f502bd;
mem[118] = 144'hf5500fa00f89f0ab0dfcfb2a00fbfa23023c;
mem[119] = 144'h060c0758f477f4f60e3e04e10215089a094f;
mem[120] = 144'h08c9f3fff717fc18f796095f07b5f2b50574;
mem[121] = 144'hf1a3f176058ef3da09b2f31a04b00989fafa;
mem[122] = 144'h041cfe46024ffba50b0bff160400fac0ff1a;
mem[123] = 144'hf416fba10ea005dcfe40fb9d0fbbfee30752;
mem[124] = 144'h089df217045bfdcd0ed30c440b1106f0f4ef;
mem[125] = 144'h0064016401440f8f0291feda0acc0f73f834;
mem[126] = 144'h0ed30f94fa9efdbdf3c309a50d9709f2fbbb;
mem[127] = 144'h0de309170b75f0ccf651fe6ff7ddf57cf731;
mem[128] = 144'hfffc045af4c3f2d3ff260c210e510285fce6;
mem[129] = 144'h03f8f875f7a709950fd4f81f061809ba0e39;
mem[130] = 144'hf89bffedfe930c8cfa38fa0d0dd7ffedf396;
mem[131] = 144'hf0270d73f571f82e087201a000a2fb05011c;
mem[132] = 144'h00700e1cf5070716fc21f198f89503aaf9cf;
mem[133] = 144'h0c15f12efdc6f4770938fef80092f81c0b3e;
mem[134] = 144'hff17f25ef13d0fa206a70f2a07e90852fb37;
mem[135] = 144'hfb3503010d360fa1fc580e3e064af68cf1aa;
mem[136] = 144'h0bd8f025080bfb75f2a2f30d05290002f3a2;
mem[137] = 144'h0ae8fa0b07ae008c0711fcd6f419ff43087e;
mem[138] = 144'h013f0f3a013eff38f10a0095f3b60fd6f705;
mem[139] = 144'hf7f904c60c4800eefb18f4d4f6dd0c34f4e1;
mem[140] = 144'hf272fba009640f8afb4b03ae0e53095c0ded;
mem[141] = 144'h088bfd3bf55b0219f1f60e1df86cf9110d00;
mem[142] = 144'h091208420ae30db106f7f1a0fc6afb5cfca5;
mem[143] = 144'hfa420f37f9300585f5c40522febc08ccf335;
mem[144] = 144'h053e0be90af5f0fef664ffc9f6d6f76ef803;
mem[145] = 144'hfab70cc4f55204b4f2f1f6170771f4590934;
mem[146] = 144'hfdcaf20906970ad3094c0481f1150dadf76f;
mem[147] = 144'h0e10fb6b057dfed20110f0aa0e20f4400051;
mem[148] = 144'hf5ebfe3bfb40fd170af4f7dc0e46f6d50ab0;
mem[149] = 144'hf4d1ffde0c6bf02009e8fed90316f00cfbfa;
mem[150] = 144'hf768fb6407b8f2980e71f3b2fcab048bf531;
mem[151] = 144'h06b0f35cf1d40b1af42f036a08070b8f0957;
mem[152] = 144'h0eabf55d08cc04c1fb3ff0f50ecb0ed60e52;
mem[153] = 144'h05b0f77ef4ad0aebf133fc1af360fdfb0985;
mem[154] = 144'h079106e0038c0c66f60dfea2f576f5aaf967;
mem[155] = 144'hf804f0e2fd51f263f799fec809e40ef904d6;
mem[156] = 144'hffd5f55cf38ff577ffb7075100e80adef48c;
mem[157] = 144'hf4d1faf209edf0ae0e6dffe701b00cd8f459;
mem[158] = 144'hff9d0e91f709fb98f1b6f166031e0f5ff9b6;
mem[159] = 144'hf02bfb60f855fcc0fae408f00c180cf9fbe8;
mem[160] = 144'hf815f7ac0d120d8ff5b40ffcfdd2fd780f7a;
mem[161] = 144'h0a4e0eb8f3600a39fe55fb49f703071cf51a;
mem[162] = 144'hfca2008a0db705a9016601c50c0d0665f441;
mem[163] = 144'h060ff39602c4fa72f22b0783f08301e3f3cf;
mem[164] = 144'h0735f38b08bd0fe8f8060e67f396081d00b2;
mem[165] = 144'hf5bbf608f8f9fd5a07250354feea088bfb4e;
mem[166] = 144'hf9b2f67502c80c970d140c9f084f0a1b03f1;
mem[167] = 144'hf6b008eaf9ff05580a30012d05c2030a0b69;
mem[168] = 144'hf766040cfde3fc9ff40c0cbb0004f402ff1b;
mem[169] = 144'hfff6fc1cfbb2056af33504660cc30d58042a;
mem[170] = 144'h0d3fff85f4e40a60f0750724f55401ca00f6;
mem[171] = 144'h09cbf72a046607b30b9afa900606fc93f19d;
mem[172] = 144'hf28ff41af347081d0ea605a7f25b0edb0d08;
mem[173] = 144'h076e07b80cc8069000c6f06c0faf0ec105d1;
mem[174] = 144'hf789f0dcf67a0bcd0e0afd35f9a4fb12f5c1;
mem[175] = 144'h0d61f45dfa7efdb8fdecf65d00720df502c6;
mem[176] = 144'hff2bf963042df43b088bff4af0ef0f600c06;
mem[177] = 144'hf9c806f5099ffc22f8d1f4ef071df5daffcb;
mem[178] = 144'h0352fa0e0a37f55ff739052800a60606fa4c;
mem[179] = 144'hf88ff7f505370802f6260a9a074bf690f4fb;
mem[180] = 144'hf13c0baffa3f03bbf921f3850bd606c9f3b2;
mem[181] = 144'h0d8d0e72f9640c65088b0e8efd0f04c4f94b;
mem[182] = 144'hffc3fcaf0e93f786f5b60afbfeb70b3e0199;
mem[183] = 144'h036b0394f741f8810b3402f1ffb6fd96f349;
mem[184] = 144'h0a0d0a15f242fffffea30765f4d80ee602f6;
mem[185] = 144'hf965f8d9f07d0d780fc001c7f858f7fdf7fd;
mem[186] = 144'h0cb50134092c0b9d01c70567094bf3b4f80f;
mem[187] = 144'hf44006d0f20506e809abf4320b2f0c8ff9c5;
mem[188] = 144'h03c1fefbfd9900e00f1f0202f050f8380db2;
mem[189] = 144'hf770f7730b11f5bcffb5f97208a50187f288;
mem[190] = 144'h02afff880ea2f806f5f100940d3bf2130db0;
mem[191] = 144'hfac4070207ce09140bb2fea30c1a04d306a5;
mem[192] = 144'h0093ff6cfb5907a4033cfbe50f59f461f690;
mem[193] = 144'h06a30d9c0f34017006bd01800de9fcfdf457;
mem[194] = 144'h08920b4cf144f79405e7f3e809baf004fb11;
mem[195] = 144'h081cf4f1fe6509a6f05a0ab9fcbbf3c1fd0f;
mem[196] = 144'hf59bf12301b6fb4b01f30ea7f381fd02f475;
mem[197] = 144'h08e608430209f4f5fa85f8d8003afc93f29c;
mem[198] = 144'h0ae9fb8cfcc809d10540f3c00c35f8d70b28;
mem[199] = 144'hff10fb400bb90cca0870f926fdeffaeaf58d;
mem[200] = 144'h0818fe5805420da5f2e5f2ebfd2309780333;
mem[201] = 144'hf96bff35f7cdfe350a7ff615f24cf4d8f00a;
mem[202] = 144'h0643f91ff4a60e42f1a00fa2f8720252f80a;
mem[203] = 144'h0be90d77fd6c089a0d6a00060f94f1a6fb40;
mem[204] = 144'hf9f305470574033bf6e30a23f3e2f06e0bd5;
mem[205] = 144'hff59f0f709bff39cfe0d0d89f2a60d720f9a;
mem[206] = 144'h0f6ff7050817f92cfbae0435f7ab005ef05e;
mem[207] = 144'h0fcdf75cf4c20d28f1190e13f44804cf0614;
mem[208] = 144'h0482f18af1fd05770d0aff4dffdcfdf2f425;
mem[209] = 144'hf22df8b2f79304ebf2eaf66ef706f92100a7;
mem[210] = 144'h0dedf01b0ec9fdabf170055ffe29013a0d7a;
mem[211] = 144'h04ed09fd093609900ee7f0f905d7087f0618;
mem[212] = 144'h0b28f724fc26f5ce0408fb0d0cbef7c6fcef;
mem[213] = 144'hf4f5035d084af9ce02830d92f4dfffc00466;
mem[214] = 144'h0a2708f100680373f2e2f4d9f896f36dfcd5;
mem[215] = 144'hfab503b10bbaf8420c40fefd0d64f169f03d;
mem[216] = 144'hfb03099ffda3fd73069b02a6fd010f09fc72;
mem[217] = 144'h0d8e0e1e0af9f5fe0b64038ef9a6f0a20af4;
mem[218] = 144'h075af5200399f8edfa840edef24d05bb07d3;
mem[219] = 144'hf9c10201fdf40a3cf754f1970481f9c3f0ba;
mem[220] = 144'hf2cdf749fed8f4e50bc8fdd503c4f2cef965;
mem[221] = 144'hf596f3dcf3c7f1360cf0f771016cf4100107;
mem[222] = 144'h0308f87efeb2fd410066f8b70ba50a7bf507;
mem[223] = 144'hf72cf14e06bc0f0e0fdf0bc7067509430e81;
mem[224] = 144'h020d0b1ffeea0d660345f3c3fd73068f0c32;
mem[225] = 144'hf05eff1b05e20914f1cbf8570a270852fc28;
mem[226] = 144'hf434f67b0c6af0cd025205c5fb16fd370c6d;
mem[227] = 144'hf9140426fe950c0d0aa10d30f256fea108fc;
mem[228] = 144'h0a8ef46a0801fa44fe640c2c045300f0f519;
mem[229] = 144'h0df9fc5c0d010ebf09c7f82af7c1039a0ddc;
mem[230] = 144'hf1d301730963f8ef0f7e081206d5037ff1ba;
mem[231] = 144'h07d5ff2e0b960b5106520387fa85fa32f923;
mem[232] = 144'hff5ff0eb0db4fd63fbc2fc00f43b0d51f2b8;
mem[233] = 144'h0f24fac40cecfd16f790fa560558f7880597;
mem[234] = 144'h070e0503fa58f18afeabfea20ab0f44ef84a;
mem[235] = 144'h04030ad7f3f20c82fd8d0a7a0ec40b66fca5;
mem[236] = 144'h0d68f63705890838f72e0cb7f1c7fc440fb5;
mem[237] = 144'h08c40a30fcdd02e4f3ddf8490d64f5a4f1da;
mem[238] = 144'hfcaa0a57f9d909760be0035df47806d1f3d5;
mem[239] = 144'hf98c0997f274015dfd100e17f7e705fff1ed;
mem[240] = 144'h008afe56fe27f6b2fda70608f775f0e40069;
mem[241] = 144'h08a90e72f789f961076ff0100a580e7ff9e9;
mem[242] = 144'hf8140c12046bf8910fb00da0083204190946;
mem[243] = 144'h012205190c9ff2cbfe3ff30908400739045d;
mem[244] = 144'hf686f9ae0f85f82d0ba9f8d5033b095b0e38;
mem[245] = 144'hf1e00cf7fb920ef5f4fe08cdf60af40f016b;
mem[246] = 144'hf49406b5fca704ba0793f59df431f4ff0ff0;
mem[247] = 144'h053a03eaf784fd52049e08160112f992f03b;
mem[248] = 144'h0eb1f0fc07e1fffd08360899f99500e3f85e;
mem[249] = 144'h0f28fcbefa72f3820faa0bbf0402099bf09e;
mem[250] = 144'h05110003062cf5150bd2f240f3ed0095f060;
mem[251] = 144'h09e00d7afc91f1c50d810067fd660b46f4b9;
mem[252] = 144'hf43305d4faf10c52fefaf9d2f751f074f942;
mem[253] = 144'hf7f3f42107d70ea4027d0307fd1a08bf080b;
mem[254] = 144'h04baf3130a7e0082f1130a6107f2f6f1f5bc;
mem[255] = 144'h0a820a660b540da209f80252f5cc068efebd;
mem[256] = 144'h00a6f0bff35500e8fbf107c6f1ff07f50512;
mem[257] = 144'h05680117f804f3adf7880a1507e80205ff88;
mem[258] = 144'hfbf0f6d6f04a0f29fb770a4cfb520133f22e;
mem[259] = 144'hf1db0538f23a053c0fab0b1ff183f35a0289;
mem[260] = 144'hff99f822fe4e0e0f0e8606dcfefd08b0f427;
mem[261] = 144'hfbf000e9f98f0b2802d5f9a1062df8d70536;
mem[262] = 144'hf7fe0098f5240c28f6a30306fac9f184f160;
mem[263] = 144'h019a0450fb74f284fdc0faff01da08770842;
mem[264] = 144'hf271fc10fb700bb8fefe0a55055e0edcf856;
mem[265] = 144'h04a1fc20f2c7f436fc220800f255f196fa86;
mem[266] = 144'hfa260e510363f3bb05d60c000a4a02e6fe76;
mem[267] = 144'hfc62f7d80231f0d0f122f62907ac0278f4ed;
mem[268] = 144'h0fb2026e09250ad60b8706d4016507c0f81a;
mem[269] = 144'hfca7068c08b9f398f937fa88f044f0f8f0dd;
mem[270] = 144'h0e72f122ff32fcbb000309de0b340ec70919;
mem[271] = 144'h0efefece02dffccf0e5e0c6af85bfecdf19d;
mem[272] = 144'hfaf4f370f98ff6460dfdfc3c0da5fdaa0282;
mem[273] = 144'hf3ca0142014cf655f7b8f36b09b8f86a0f84;
mem[274] = 144'h0f93f9ed0f15f9d601a5f57e0191f6e4fd56;
mem[275] = 144'h057b017e043bfff9095b00b20454fe010ef5;
mem[276] = 144'h01210765f2580c880a1bf1910070fbeff748;
mem[277] = 144'h060907f8032f0c730e08f82e01430a790d47;
mem[278] = 144'h0c5d02790208fbf4037dfea400a5fbc8f401;
mem[279] = 144'h07080c2afff50db3ff9d0ddcfae90ec40c0f;
mem[280] = 144'h0562f995fbe50d9d01dd0b26f323f830ffe5;
mem[281] = 144'hf4aefa9b035df39d04ed07fffbb70c490875;
mem[282] = 144'h003f0419fb580611f731f65902b8f47bf6ef;
mem[283] = 144'h061ef0f001dbf2b7feb1045b0f72f7870cc2;
mem[284] = 144'h0ac9089ff735f9980cacf71fffc9fc180039;
mem[285] = 144'hf67b04bef13ff8670859fee00d84f0ef0daf;
mem[286] = 144'hf3d2f5ee0cf501a8f7b3040d06980a23f1be;
mem[287] = 144'hff4d019606dbf442f11407670e610556f6c1;
mem[288] = 144'h0c540bde00b9f2050fae0722082f09e70c61;
mem[289] = 144'h086efca3f6e80fb00681f5360db10f5df235;
mem[290] = 144'hfacafaf0fc5502310da00e4d0c5701a6fc96;
mem[291] = 144'h0d7cf92509c8faa9ff9ff07dffec01cd00db;
mem[292] = 144'hf6410467f3360f9d070af36e016efdf3f0db;
mem[293] = 144'hf0ccfcf4ff80fac9fdd0f48ff33e0ba60237;
mem[294] = 144'hf7f3f709031b0bb1fa9b08f8fa940dcffea8;
mem[295] = 144'h0dcff24601870a3ffefbf4770ed9f310095e;
mem[296] = 144'hfc92fa1cf4dffe8af8d1feda0d060018f6af;
mem[297] = 144'hf60e029df6c809750b70012a0d62fbda006a;
mem[298] = 144'hfddb0c33f4e8f079ff7e0eb6ffee0d360b49;
mem[299] = 144'h05290704f99607acfd93f04ff50901dd07c9;
mem[300] = 144'h05e7fc3cfa9afa6304d9f54904e7ffd8fbee;
mem[301] = 144'hf7dcfad30ba2ff9befda00d3ff01f2110cea;
mem[302] = 144'h0ccc056c0d37f10a08bafcccf3c1f8affa54;
mem[303] = 144'h0c4af92af3d4f116fcd4074d0e7df0eb05d4;
mem[304] = 144'h07f00de1f79d0a19f62f0b4405a8095b0aee;
mem[305] = 144'hf30ef5c2fc8e03c8f7760267f29200aef5f2;
mem[306] = 144'h0cab0999fcb4036ef84ff65f0ada0b65fcfa;
mem[307] = 144'hfedcf314fa0b02a3f401f40400c70b60f93a;
mem[308] = 144'h0d410f35fac20e4af3c90b7c06160f920c81;
mem[309] = 144'h0c4afa76f78f0bcdf84e0fa4fb4cf1a90d30;
mem[310] = 144'hfbcf05cc0a440d260440088e0604f67f09ac;
mem[311] = 144'hf83c048fff4f0db50295fb32ffda0e3df848;
mem[312] = 144'hfc5df72205330499f4cafdee0bf6ff5dfb21;
mem[313] = 144'h0e02ffeffecd0d45fcf4010909e9f61cf065;
mem[314] = 144'hf1f10ae5f80b097004d10d9cf32903bb0461;
mem[315] = 144'h0363f14ff77d0a140f08ff60f4220ea10045;
mem[316] = 144'h0da8eff1f467f4bd0c26f53d0f4a0ca10b88;
mem[317] = 144'hf0eb0881f487f79e0f22f4880e5102b1fb2c;
mem[318] = 144'h0209037a0e6bfe6204bffe22fade016ef7ba;
mem[319] = 144'hf5c2016704cffa16f342fc660ea60a42f1ce;
mem[320] = 144'h075ef3cff21afe460f9f0caf09aefe65f7c4;
mem[321] = 144'hfe3cf442ffd90783032300b10d4c00e20bce;
mem[322] = 144'hf75d020f002e0ca30a68f6bdf792eff20ef2;
mem[323] = 144'hfb910a780112fb19f6aa02c107720d25f61a;
mem[324] = 144'hf90bfa98f94d0bf0f28ffd7202040cad0709;
mem[325] = 144'h0d2f07b30bb8f87e0d9ff1ac0bf3ff6b0d70;
mem[326] = 144'hf9a4fa750f910ceb004201ae0b3ffd83fcbb;
mem[327] = 144'hf5cf03b10aaf042406cd01670bec0bd903e2;
mem[328] = 144'h0f6e0c20f5b6086ff6c903bbf35fffa5f638;
mem[329] = 144'hf7e0010e09e8fe110201f263f842f9affa26;
mem[330] = 144'h07d4fb20fed8f7e5f662fc44f31b07b1f433;
mem[331] = 144'hfdf0018dfdb0f5c50685face08be02d10e32;
mem[332] = 144'h0217f33706f8f29f06b100f3f0bdfe17f234;
mem[333] = 144'hf11d06dcfb3af6adfece0871f4b60744f92d;
mem[334] = 144'hf7a3fff80c5406faf3e7f89404cc032f097e;
mem[335] = 144'h0bb00bf50a25ff37096a0a8efa8eff37f8da;
mem[336] = 144'hfdc102660ec409cb0e1af80bf5e5fd1efba7;
mem[337] = 144'h05b6f7aaf0200b9cf2d108860d9bfdfb0f70;
mem[338] = 144'hf6f50a0001a6fcabf591f038fdd6f3f1f79c;
mem[339] = 144'h0d4dfa0e0bb6f69a0a850704f8c4fb34f6e4;
mem[340] = 144'h0e6efd760d57f5300ad80200f6860788f687;
mem[341] = 144'hfde109ac01000944f5aa07cdf3880a71f92e;
mem[342] = 144'hfd98060ffaf10c2309200bb00d2c001c0822;
mem[343] = 144'hf891fdc4f6570f8700ae0e35ff9c01f1f1af;
mem[344] = 144'h007dff930c3efb2605570d0405ddfa4c004d;
mem[345] = 144'hf6fef605f0bffb480050fae9fc80f33bfead;
mem[346] = 144'hf257082bf76e0d170f46f0d9ff6308cf0946;
mem[347] = 144'h0f41f1c201230aa20d3cf5fd06f30e2b0721;
mem[348] = 144'hf91bf2f10864f37ff79307a2f1b7fa3607f1;
mem[349] = 144'hf309f28d0a44ffacf2c205e8f2e3019b0d57;
mem[350] = 144'hfd04077ff4e70c9ef8e40c35f405f720f1cc;
mem[351] = 144'hf807fec7f239f886f0a5fcfff19b00f9fcb2;
mem[352] = 144'h0b65f9480625fe16f87e018f05d90d980041;
mem[353] = 144'h0951059d078f050d0cd604430712fa4fff82;
mem[354] = 144'h0fb5f2bf0ea006220c27f99d0a8308c9f36e;
mem[355] = 144'hf05703290116f858fa58f12ff79dfbe9fe01;
mem[356] = 144'h05dcff5f0027f4adfb370772fc01f710fae6;
mem[357] = 144'hf74bfc85074f01e10fb4f9b00bd20d640e19;
mem[358] = 144'hf4120f34f005f6e50015f7130bdaf664fadf;
mem[359] = 144'hf4b7f681f4560411f99a05ba06d4f49f0781;
mem[360] = 144'h04fff120f04a0437f82208a9fe7d062f05ff;
mem[361] = 144'h09fd0d770f9507eef845062f05b6f6cc01ad;
mem[362] = 144'hf526fd70f1b5f8850d7004ec0bd4fe6e0236;
mem[363] = 144'h048c0ca30290f138033f0113f7050226f540;
mem[364] = 144'h0361083400930a890f47f5920eeff23df181;
mem[365] = 144'hfd000985f54df19108100bfcf6bdfedff2ae;
mem[366] = 144'hf14a04bbfc15ff7a0cf6f838fa5803410d23;
mem[367] = 144'hfece0b8702a001610557f417094101c20a5e;
mem[368] = 144'hf149f28f0558fa99f3560521f7c901890c61;
mem[369] = 144'hf87b01b4038bf09c0042f96bf47f000307c5;
mem[370] = 144'h0e67f6180b36f679f8f2f8c7f4e2f0a7098a;
mem[371] = 144'h0dafff000965f32707a2f5a30850f3450224;
mem[372] = 144'h03c50d1d028904cb0cfa0ebf042ff2360314;
mem[373] = 144'h037e08cbfcdcf1fc06f805e906d609a20a0d;
mem[374] = 144'h08cd068cf204f05ff53d09de08a603fffb01;
mem[375] = 144'hf542045ff0f5fdaefcdaf706fc220717fab7;
mem[376] = 144'hf3e806aff1cef552f33a0be10afff8d9fe68;
mem[377] = 144'hfe1a0854fd96ff670a72f8caf029fa8f0028;
mem[378] = 144'h0a070c7a00aa0e7af3b1095af300f1eaf3e2;
mem[379] = 144'hf01400b803f3fe830825f6d1f72ef5cdf5e8;
mem[380] = 144'hfebd094504960503f8770787fa9f0d7ef78c;
mem[381] = 144'hf350f1a409d407eb01910a3efd29fafb0a17;
mem[382] = 144'hf19b08080f47fb970dadfa5204ff0ae9018f;
mem[383] = 144'h0a17f1e3f7c7fe77ff700d88f343fa230182;
mem[384] = 144'h00cc0ed4f0920e79fc7e0639fcdff2f2f196;
mem[385] = 144'hf1b3fbaafac508900400086cfa8ef5170845;
mem[386] = 144'h045703fcff0ff1fa0b2e02c30841f48df13a;
mem[387] = 144'h05ff05100294f4bbf514f7700e8805090d4b;
mem[388] = 144'h018f024ef1a70945027ef1e4007cf2d50399;
mem[389] = 144'h0dca002c06e5037b00ec049ff5790f7b00bd;
mem[390] = 144'hf6a80326fee9f2ec0030f49d07e9f0660396;
mem[391] = 144'h0981f19408e2f8d7fac5050d0c78f2dc059a;
mem[392] = 144'h03ef0462086af8b0056bf54ef642feb00eb2;
mem[393] = 144'h084a0c18fe8d0223fe61f49cfe2a04430523;
mem[394] = 144'h0af4f70c0d37fb430e080e9f0627fa750272;
mem[395] = 144'hf2ab06fd06adfbe0fb31f0c20251059cf652;
mem[396] = 144'hf77bff510d34071ef21c04fb013508f10eaa;
mem[397] = 144'hff87fd21043700a40c58fdd4f27dffe1fd09;
mem[398] = 144'h07a506f20fa1076e00c6f3d3feacfea6f0c7;
mem[399] = 144'h064e0649fc16097602d9ff9cf3b4032af972;
mem[400] = 144'hfe8007aa02c00f0f055c0ec0f3f60726f9b7;
mem[401] = 144'h095ffc46fc96073c0583f6ed04b6f0760497;
mem[402] = 144'hfffcf1fa0c0f03ae09b7fca00bd8fa020e79;
mem[403] = 144'h0a3ef84c0bf9fa14075f06b1f516f6fbf9e2;
mem[404] = 144'h08e4fd98f884f21ff19bf3d3f41ff865f218;
mem[405] = 144'h03fcfc330643080df8b0f3b30c4601e409eb;
mem[406] = 144'h092af5550f8e06c90a2a025e064c09ef0e14;
mem[407] = 144'hf6e906be09660a4af85f059f07770070fa2b;
mem[408] = 144'hf3280e43f179f6c9f5d50c6c051105c70825;
mem[409] = 144'hf4bbfed40553f5bdfc30036bf2c5033d01ea;
mem[410] = 144'hf73f022efe880926fcf8019ff417f099f8d6;
mem[411] = 144'hf6aef43affe1fd6b06cbf81ff0e5ff02f111;
mem[412] = 144'h0a53fadf06810438fb6909fc0c76f6550d0b;
mem[413] = 144'hfba80a93f456fcc9f847f41cf39af8c3f796;
mem[414] = 144'h0583f1e3f739039ff0ccf09001ad017d0aae;
mem[415] = 144'hfde402da0ced06c0f710fd1b0c8500f403f4;
mem[416] = 144'h0abdf429fcb9fd3cfbf3fd440277fab80035;
mem[417] = 144'hf7d801c2023e01bbf8df0beff2ce0298013b;
mem[418] = 144'hfb7507c6fc790604f60df5f700110cf309a7;
mem[419] = 144'h0b72f91afe2e0305f1b708a8fc1d0bb9f8fe;
mem[420] = 144'hf776fe8a090df7d3f6e6f42f0a8df4d8f5a6;
mem[421] = 144'hf1c1fc40f9840ea1f403fdf0f278f20a064a;
mem[422] = 144'h0b490afaf143f9defdb8fc470327facff5ab;
mem[423] = 144'hf223061804e70dbefe0af2360bc6f095f6d6;
mem[424] = 144'hf130052d0c0afd41fbabfd210133f66ff06d;
mem[425] = 144'hf2f002b3f9f8fcfe0939018600b3fa1906cf;
mem[426] = 144'hf425f46aff04f304f79504f2068d02040dbf;
mem[427] = 144'h0d32f860f8dcf305f5e00b7bffb2f3c30de1;
mem[428] = 144'hf8f507b8f86efec9fa740e290a68068803f8;
mem[429] = 144'hf7f80f3d020f02a90d6b041bf5b0026bf289;
mem[430] = 144'h06560e03f6f00da5f6bff564f76205d0fe67;
mem[431] = 144'hf1a70a9e0108f6420a9df340faf70437f001;
mem[432] = 144'h0c5ef93d0c0c0fcc08520862f5a00a59051d;
mem[433] = 144'hf732fa6905870afbfb5df4ea0474f8c3fc3e;
mem[434] = 144'h08650339f188f97f0f37fc76021e03880eab;
mem[435] = 144'hf37d0605f2f7f4e706bb02c2f314fc7c03cc;
mem[436] = 144'hf3ba0e700130f04df49e09a80adcfba7f585;
mem[437] = 144'h0f840c14f282f236f431f8c5064cf2890bec;
mem[438] = 144'hf028ffabfba4f6b6f4df04ac0586f5a8f3b0;
mem[439] = 144'hf635f1e206230e85f31bf33ff7c2f3b80531;
mem[440] = 144'h0185f8e60898f90b0141044dff7901260cd7;
mem[441] = 144'hf576fef3fcb1fbd9fb4bf2ecfc69f2430f0b;
mem[442] = 144'hf28cf308fc6a054bf0c0f6fafea1f9a7fbd1;
mem[443] = 144'h068df7f2fb95ffb50e74f84df7440cedf2f1;
mem[444] = 144'h0bc4f381f2edf63efa0cf346f958f6a90f43;
mem[445] = 144'hf7a8051f02f90b92f8600c8d0f4ff4bbf311;
mem[446] = 144'h037cf725040bfb98fecaf699fa6ef98a00af;
mem[447] = 144'hfab009490dfd064cff5af83efe17f85af09a;
mem[448] = 144'h0cc50484ff22fc34fdeaf2b7fbdefcb806a9;
mem[449] = 144'hfc64f4d0035c0697f4400550038b033403bc;
mem[450] = 144'h08e00959f9cb0249f7e7f4c80b03f07c086d;
mem[451] = 144'h067f0f230db7f200f3c60bd90de3fe82f703;
mem[452] = 144'hfb4f02a70e12f770fd52f520fa5905cb0b68;
mem[453] = 144'hf93d074803b6f6f107c2f3ec05300f0401ef;
mem[454] = 144'h0a4ef833f560f391055c0146f969f8a0fea8;
mem[455] = 144'h0d1f03e7f153f552f466ffe40da0f308eff8;
mem[456] = 144'hf52c08d0f31afe6ef305f388f97bfc30006f;
mem[457] = 144'hf678077a094df329f21205dd0f8100240d3f;
mem[458] = 144'hf645fe080f68f8a00366ffcb002afe0af0e3;
mem[459] = 144'hfaef0938f9b3fe6106ed0678f30909090eaa;
mem[460] = 144'hf32ffb740201f2ebf7e20757039a06200eec;
mem[461] = 144'h0ab9ff400edcf0f30f48087c03b309d0f2e9;
mem[462] = 144'hfdb506f0f4f70af40a3b0a7b0bee0db70747;
mem[463] = 144'hf418f766086ff54601b0fa48f0840fb6fbf6;
mem[464] = 144'hfed3030cfb970bb4023c026a00f20ca70450;
mem[465] = 144'hf0490f0cff240f1d0124f883f99404fb0a3d;
mem[466] = 144'hf0ccf4fbfa18f9f108bb0a820f5bf9df0354;
mem[467] = 144'h0179f901fd48f0100f4efe870991f5ccf576;
mem[468] = 144'hf330fc860134f8100bf100d1f511f344028b;
mem[469] = 144'hf793086afed007e3fabb013605ecfe450594;
mem[470] = 144'hf90ff6830bbbfb82f8a6fc2e0142059c0f3d;
mem[471] = 144'hf96c08dd0dc2f5a70b58032bf0bdf47507ea;
mem[472] = 144'h0923f22bfe1707d7013e0af60e3e095503f3;
mem[473] = 144'h00c4f8cf064a0da4f791f9ce04f60170fc15;
mem[474] = 144'hf9f4059cf1c009af0d2103e30c1b00460cfd;
mem[475] = 144'hf8120c6f002f06f3fc9f078a0d0f0140efe3;
mem[476] = 144'hf4b40a8901b5fa35f17903750cbef048f2cb;
mem[477] = 144'hf04407a7fdb6094cf2840c7efabd0d1afc2d;
mem[478] = 144'hfa7a0ba8fb970099fa8d009e08f70bb8f2cd;
mem[479] = 144'hf1690515056c0ff4fb540f150915f3ea0abd;
mem[480] = 144'h07a7057b077ef4f6f9d2f2e7ffaeff51ff7b;
mem[481] = 144'hf631006f0a9103a4f75af269f172f67a09be;
mem[482] = 144'hf1a50766fe8b09e509eaf4bb0943f6230fa1;
mem[483] = 144'h00940b3b00d708c402f70f610752f217f081;
mem[484] = 144'hfc2f01dbfd2d0d2af2ef06700b6e0c62f669;
mem[485] = 144'hfc5bffc20e7c0576fbdbfa7d0f4e0c9ef0e9;
mem[486] = 144'hf35e0d53043afaa4fbecf4a40d9dfe4e092b;
mem[487] = 144'h007ffe4402fc0e51020bf2440900fa510794;
mem[488] = 144'hf439f9370276f74900720d14f25bf5280709;
mem[489] = 144'hf7f4f40b07a5081601e70d57027407a7f942;
mem[490] = 144'hf0abfd1509270c5704a9fb19f1170c58f550;
mem[491] = 144'h0908ff16f659fd8b0829fa0c021907c50363;
mem[492] = 144'h06d40eca0342f833f110fa170c6f0aaaf0db;
mem[493] = 144'h0f6ef9ac04bff870f31c0f340afff2b3f123;
mem[494] = 144'h09adf678022f0be709a3f53efd170355f136;
mem[495] = 144'h062606270d9ef9eaf9c00ec0050af3c401bd;
mem[496] = 144'hf6020a050f85fb2e011e06510e15f8c6f56e;
mem[497] = 144'hfbd30827fcef09e700df07a6f7ca0eb00501;
mem[498] = 144'hfa41081dff87fbb0ffd605b9fb23f8c701fc;
mem[499] = 144'hf9fe0cd0061b05d3f894f84e095d09030084;
mem[500] = 144'h0f4b0f910ed9fbc20dbf0fb1fa28fef3059d;
mem[501] = 144'hf837fcfafa9a0223fd0df1e1f1b90d230844;
mem[502] = 144'hfd5c08ba0c570375fc89f70a06930cadf503;
mem[503] = 144'h0f64f4edf4580438f32d03c6f4df09960196;
mem[504] = 144'h08f0fa830352f21c03a1f4d9fac7054bf0ac;
mem[505] = 144'h0f290c0b0240f2e2f32808ef084f0ddef8aa;
mem[506] = 144'h0874fa4dfc16f0ba040c02880b43f386fd65;
mem[507] = 144'hfa450318f2a70602f4770746f3620d780ecc;
mem[508] = 144'hf1bcfd1df502f690f78b0914f2760a1ef16a;
mem[509] = 144'hf2f507caf70d01eb04f7f74d0bbcff07f6f4;
mem[510] = 144'h0bd8fa25f62cff55f6b5060ffb33f23ffb0b;
mem[511] = 144'h08a4f324fa24ff05f721f072f070ff3cf04e;
mem[512] = 144'hf4b70b40ff95fd3c0a500ad2fa220523f47e;
mem[513] = 144'h0326f397fc55060f0ef4f2aaf1b1fe46f620;
mem[514] = 144'h09650c25069006510d4907cafff8f09dffa5;
mem[515] = 144'hf5070a95f1abf3bffd9805df024c0985f00f;
mem[516] = 144'h03a609130322f0fe0dd80350f8a0011df324;
mem[517] = 144'hf6ed0b9e05f7f4920aa0f2d103910e90f593;
mem[518] = 144'hf4e609650846f045f435f9d20871f90f0913;
mem[519] = 144'h007e0d820872016c0413f8f9f2220efe0fb1;
mem[520] = 144'hfd1ff66cf690f226f50af4a6003efa0f055e;
mem[521] = 144'hf142f79103d4facf01c600fd0952eff108b0;
mem[522] = 144'hf88b0f000336051bf6f8f4dafc070662fb2f;
mem[523] = 144'h0742fdd0091900b3f2e2fe32050c050b0603;
mem[524] = 144'hf06b00f10fc1fda6074df1ff03b50a910552;
mem[525] = 144'h0f2cf973035a08fa0bb50f0a0af506b50b43;
mem[526] = 144'h0905f97609bbfb5e086cf6820cc303f50fe5;
mem[527] = 144'h0371f6960bfdfdb902f5f03bfe060df308c1;
mem[528] = 144'h073ff51bf3cf06e3f42c09a8f20703c00e14;
mem[529] = 144'h07f004e20dec0f25f007feaaf745f2a7fec7;
mem[530] = 144'h0424fdb4fbbd0442f331f069f8230a91f816;
mem[531] = 144'hfa38080bfae207000dc10314fb90fec401c6;
mem[532] = 144'h026df2d20e1d04cef879f9540b8af298f021;
mem[533] = 144'hfbc1f7e9fedc0f0403c5fd02ff5908ce01de;
mem[534] = 144'hf1c1f40bff72f2d00edbf354026901d606ed;
mem[535] = 144'h02200e6f03b004aeff5ff1330b56fbbefc35;
mem[536] = 144'hfa1402bff4e6f7aff8aa07310feefabb085b;
mem[537] = 144'h09100a6af65cf873f444fcdd0d14f529fc66;
mem[538] = 144'hf9610562019506f901a8f284f433f57b0047;
mem[539] = 144'h0481ff2fffcdf1a1f63109b2f734ffc60e15;
mem[540] = 144'hfa41f0fefb0e09110749fa3c0d9f081f0a72;
mem[541] = 144'h01eafb26f576f4eff76bf4d0f8bc0e090f7b;
mem[542] = 144'h0d80f143f825f1e3f3880385078ef3d20d40;
mem[543] = 144'hfc8afcb0f8b0faa906370076f454f4420c06;
mem[544] = 144'h0a86072d004102050505fc9e0ca50525f3a7;
mem[545] = 144'hf52d02cf0c7cf2bffea502d205a80df3f588;
mem[546] = 144'h0f45f5e50e0f0eaef42df45800190851f623;
mem[547] = 144'h0569f8400955f5090030f8d5f5050b3b01b1;
mem[548] = 144'hfe64fc1c085a0a18f12401a009a3f46f01f9;
mem[549] = 144'hf55df053f7e60f94f53d0732f9950e1c00d3;
mem[550] = 144'h0845fa94f22c018a0e8bfb2a0e98f978f9c6;
mem[551] = 144'hf6f0fc30026f0f750b24fdb901230cf20b3d;
mem[552] = 144'hfc6001c3002809be092e0130f4f3ffa5f40c;
mem[553] = 144'h06c3fd990cb1ff2607bb098af9aa0d210b30;
mem[554] = 144'hf8ccf7da0103fd98fecf02970521f8a9f0cc;
mem[555] = 144'h00aef4da01b5fed3fe6205a40fd7f492ffbf;
mem[556] = 144'h0597eff4fde9fb9609edf0a306830956fa42;
mem[557] = 144'h0de8f8a40e6e09c901a70d0802f6f4fbfd71;
mem[558] = 144'h0ab30afb0d40f3dbff5802a90b9dfe15f20f;
mem[559] = 144'hfbf00c69fe75f8f80718f93df582f24a0834;
mem[560] = 144'h0f1b087ff581fafc080cfb1b03ed05370af5;
mem[561] = 144'hfc250321017b0f88076bfd48f9c10efdffca;
mem[562] = 144'hf510f9b2f894f66c0b77f0fbf2840713ffc4;
mem[563] = 144'h00c40e4ef035f3d8f20df8ef0c5d0405f25c;
mem[564] = 144'hfe43089ff38cf2aefeed014df866f106fb68;
mem[565] = 144'h0894f31eff44f9b5f2e10b07f4ab05bbf9ba;
mem[566] = 144'h0b8cfad900920efbf072fbf2f0fb0e3df498;
mem[567] = 144'hfbdc0bdb00390a040d7bf54c009c04800e9a;
mem[568] = 144'h0ccff027ff7b0dcdfdf4f419f57b03a005e4;
mem[569] = 144'h07a8fd32f322ffcc03b1f566f557f2ac0b41;
mem[570] = 144'h01c20560f9eef5da02b9fb9af8c406f6f714;
mem[571] = 144'hf8a6f96cfc990eb9f661ffca0363f7ae0351;
mem[572] = 144'h0a7906aa05f3f608056bff14fe83fc87fef7;
mem[573] = 144'hf4e4f7f70eff05d60fdaf9baffc9f4670f51;
mem[574] = 144'hfe37f2670c7a0a26016cf188090f06aef66f;
mem[575] = 144'hf2840892018e0466fa77f8c6ff4c0edef8a9;
mem[576] = 144'hf8860c41f2d7f95000d905f90f83f72b0129;
mem[577] = 144'hf1860b8202b2f61b0c75f4a0f1130808f64a;
mem[578] = 144'h0387fa1e07b80314f07b09a8f1960a17068a;
mem[579] = 144'h03730b16f1a805ac04fb05b00cd2f5c6fcb0;
mem[580] = 144'hfd09f661f91ff04b02b30cd10cc3f8bffdd2;
mem[581] = 144'h027309a40363f197f7abfce80e5c06a00640;
mem[582] = 144'h091df71cfcf40845001ff8fe00ad08300fb8;
mem[583] = 144'hfff707740a970d07fa36f68cf44df288f5dd;
mem[584] = 144'h050605ecf3effaeef4170a7af4daf93c06ac;
mem[585] = 144'hfd410c3af9670d3b078b07880b25fb1af760;
mem[586] = 144'hff52f64f0c66083d00a3f69efd21f50305df;
mem[587] = 144'hfead02d20f6905610942f7cc00b10ef207ec;
mem[588] = 144'hf5eef569058506b30dbd055b0a240c12f2f4;
mem[589] = 144'h009908a6f602ff39f7a40c2c07b5fd0f0349;
mem[590] = 144'hfc1cf9080b1d037cff3bfdad03d1f544f5ce;
mem[591] = 144'h03fe066ef25eff7a07e5f22b0cb00ea70e36;
mem[592] = 144'hfcf80bd30cdfff5cf5b7f712045ef58efff5;
mem[593] = 144'h07a2f3e20d5a01360c48f75e07fe077e0173;
mem[594] = 144'hf9dafe270cf3f29d072bf16f044708750f86;
mem[595] = 144'h084a0af4f8bcf46efe2f09f70847f0f608b3;
mem[596] = 144'h0cc1fb4cf6cdfb810719f245f4070856f8c5;
mem[597] = 144'hfa410f53fe420ea4f2e9065c0ee0f4400e75;
mem[598] = 144'hf95a0fb3029dfb27f62a0e00f85d026f08bd;
mem[599] = 144'hfeaa0ebffaba01e40e5705a8f24600abf8c5;
mem[600] = 144'h0a04f97af977fda2f8aa00faf8eff187072d;
mem[601] = 144'h008ff9cd0c83f50bf510f8f7f8e7f8a8f913;
mem[602] = 144'h0809fde8f603f4e407b5f245fda8061f05ef;
mem[603] = 144'h0ffa09d006610af201f80ece0d0d0cc1ffa3;
mem[604] = 144'h0d9b0517f8cc0a7702c3f70af4b40b51f4e1;
mem[605] = 144'h02a0f743f44af0f7f8c6f2c0f739f06c05bc;
mem[606] = 144'hf657f147f9a20d85f4030b1cf1670a9e0e49;
mem[607] = 144'hf861fcfcf9adfe3ff1bcf26405f6f5a0f103;
mem[608] = 144'h0fa90e7af8640b82f186f5120de5046f011b;
mem[609] = 144'h038b076dfbed0a0c03e5ffa5f4d1fbebfa2f;
mem[610] = 144'hf286fb580283015b0a0f053303a2f3d5faae;
mem[611] = 144'hf52708abfb67f1d3f4a4f264fb57f3eb0242;
mem[612] = 144'hfd52f6f7fd42fd32fa9d0f3f0b680e0a002c;
mem[613] = 144'h0ca6ffcdf28ffdaff57bfda20bcef2c00144;
mem[614] = 144'h0ba1f7470ed50d2a0b330f40f62bfdb70033;
mem[615] = 144'h0d740a750be8f9e5076604dcf676f401f598;
mem[616] = 144'h0b76ffc4f41fff9804e9097e0752096e0a68;
mem[617] = 144'hfd9607dc08a50ad6f5e7f7b0f605f62ff4c1;
mem[618] = 144'h0e5e0adcf645fca603adff07099bf6f40013;
mem[619] = 144'h0f480da7f8780a12f04dfddaf46d06e0f0ba;
mem[620] = 144'h0021075af4830f710a240badf8f9029106b2;
mem[621] = 144'hf00e0477ffae0c0af8fc0a350a5cfa560be6;
mem[622] = 144'h00110c9cf85d0571f23efd7b0fd20969f48e;
mem[623] = 144'hf69cf264f466f7ae009f0b76f2c6efe9f5ac;
mem[624] = 144'hf4a9f71df8bf0c6bfd7bf8800cd5f0590f71;
mem[625] = 144'h0f9e0f9502b70d3d05380e710d540eb0faac;
mem[626] = 144'h0bf803df0cda0ae2f382fe71f27afc4ef6fc;
mem[627] = 144'hffa2ff2708fcf426089dfbd1ffc5f9e3fcdc;
mem[628] = 144'h05c3f01b000dfd4ff1de0cfb0a64f07df86a;
mem[629] = 144'h0ca4fda90ef1f6e1f5acf69f07eff3aaf830;
mem[630] = 144'h076ef8af0ecd0e290b170d4cf59109c7fc1a;
mem[631] = 144'h06e7fcb2f9b2fe06f2ae0120fb03f16b0db9;
mem[632] = 144'h0cd6fcbef1750bbfffe0f27e0556f64902ff;
mem[633] = 144'hf5a60a46f56708880ddff851fd47fb500f3b;
mem[634] = 144'hf3b7f01b07480c2b023006fd06c10167f099;
mem[635] = 144'h057d02b3efed07e806cdfcef0119f5f3f1e4;
mem[636] = 144'h04bef718f0fe09e3043dfb720776f9c401e2;
mem[637] = 144'h04870c2efe560064f152f9d8ff4afab9f3a4;
mem[638] = 144'hf1b4f64df09bf0aa0a7bf75af30703e9f2ad;
mem[639] = 144'hfe65f5ecf4c0fbb0f2e80941032af9bff978;
mem[640] = 144'h09bd07ef00c600fef8daf98b046e0db8fa6d;
mem[641] = 144'h09a1f4e501a1fedf0846f389fb40fcd9ff1b;
mem[642] = 144'h02c60dcdf1bcf142ff6709760343f0defb09;
mem[643] = 144'h08660b29f608f07200d309c604ff0741008b;
mem[644] = 144'hf126f61e0adefeca0c6e0dd2fe86f20ef028;
mem[645] = 144'hfdac064bf655f9f4f95506a4fbd2fbaff06c;
mem[646] = 144'hf1dcfb0e0fb9fa7a0222f847f5df03acf84e;
mem[647] = 144'h0558000705c4f870fb74ff710208f71405b2;
mem[648] = 144'h0e020401fc3105a8fc32f6e6f502fde40f2b;
mem[649] = 144'h01a400170d650137f886fbacf31ef9220a92;
mem[650] = 144'h092e02f7f4f30cacfa54f7acf3d90fe60697;
mem[651] = 144'h0d270c0a04f60a36f695f9c10170f8150c33;
mem[652] = 144'hf9bbfa060b9d01960c5104f9fd0f0202081a;
mem[653] = 144'h0c880851f155f796091003e50acf0cb6f7b3;
mem[654] = 144'h07090d9601130225073a04be078d0d36f2c2;
mem[655] = 144'hfa6603200ff3f53bf57bfb59fa6ff53af73a;
mem[656] = 144'h051009d3f27a0ec3f9750b50fe93fd75fa34;
mem[657] = 144'h0b70ff3d0e070447046d0087078ef356f117;
mem[658] = 144'hf97af8f7019efa4ffb07fb570143efd3f2b5;
mem[659] = 144'hf9670da7fcc9f5d9f2cd0e7df904089ffc60;
mem[660] = 144'hf5b1fe6808f2fec60a86057ff40d055a0d99;
mem[661] = 144'hf219f6b9f2a40db103dffcf103c50ebf0804;
mem[662] = 144'h051ffb9c006ef7daf9edf232f93cfb580305;
mem[663] = 144'hf50c0475f021f456fd66f08a0a81f6a0fad7;
mem[664] = 144'h049e04a8077affa7fbb10b3ff0c7fc0d0cc0;
mem[665] = 144'hf926f9fa0abbf46c0bae0c8cf01bf2a6030d;
mem[666] = 144'hf0ff0dcc08b7ff890253f5dd086bf881f2e6;
mem[667] = 144'h0ef1f90dff2205d4f395fb5ffa080006fb4f;
mem[668] = 144'h00faf8fafb25f00b081f0433fccd067b0c18;
mem[669] = 144'h01dc0baefd02f0def32dfec6f01af8900b2e;
mem[670] = 144'hf8730c97f45f0a70ff48f23efaf50c84fd87;
mem[671] = 144'h0f0d01f603690e7805a0f18206b0fe06f5c0;
mem[672] = 144'hf629fe1402350cc6fe2af655f91bf2b0f7e8;
mem[673] = 144'h0599fce40d4ff90fff58f7180ee9fc16fddd;
mem[674] = 144'hf560f7d3f01806b208c3f0cf0b63f0390436;
mem[675] = 144'h0ad7f0c60634f2440cd00fccf493f4c1f225;
mem[676] = 144'hf30105d102ad018afbef073ff2a10202ffd2;
mem[677] = 144'h04a3f27001600f21086f0d5706bafb98f040;
mem[678] = 144'hf252014e071afe5bfc60fac3fc14f1dff373;
mem[679] = 144'hf48508c4fac9088b0f8b0c380e560249ff62;
mem[680] = 144'hfc45f20f04fc0b9e0bd804020dad0147f1f1;
mem[681] = 144'hf84009fef62e033d03da0b2af15af3fbfd29;
mem[682] = 144'h0f5cf92ef104fb30f185f1a800cb0f37f717;
mem[683] = 144'h0bcffde30c76f27dffbb00a5fa150541fbe7;
mem[684] = 144'h0e16fd100d95f399093cf4540d34fcd501a4;
mem[685] = 144'h0151fd650e3a0e6c0ac40cc2f3d9fa55fa9b;
mem[686] = 144'h03e20fe70dabf63cf224f4bef1f20bcbf6bc;
mem[687] = 144'h04f8f898f1e409cb0b52fb0100c4f18efd49;
mem[688] = 144'h054902e8fc84fbf7f942f0ef0cc3f2110deb;
mem[689] = 144'hf6080d9204b8f101f5590e6d0169fdebf068;
mem[690] = 144'hfaa60d3af4aa0b5df8faf6c30468f521fbf7;
mem[691] = 144'h0584071c0a7ef1270bc4fd67f9a4094a08ce;
mem[692] = 144'hf3f7fefa009001030876f2c0f592f791f707;
mem[693] = 144'h0aa6fe90f517f2c300250448f1710d89f85f;
mem[694] = 144'hf2dd015af4700773083a0c0f041007b905a4;
mem[695] = 144'hfaa30cfcfe7c034208c1fa070132fda7ffbf;
mem[696] = 144'h0dbc03d40e97ff38045b06740799fc750811;
mem[697] = 144'h02f90b93fead0cd1f243005c024afef6f582;
mem[698] = 144'hfffe0a5dfd5cfae3f4b5fdbd078106bc00f1;
mem[699] = 144'hf109ff01f2a8f693fc1ff35c08290501f3ef;
mem[700] = 144'h0778f294017cf129fc35f68007e4f5cf0df5;
mem[701] = 144'h0c06f83afa5bf36208b50b59feb902850740;
mem[702] = 144'hff4e0b1dfa79f7240176f036f770f184018a;
mem[703] = 144'h0014f7730e73fe980718f5fc02550f50f396;
mem[704] = 144'h0913fe5dfa40f4f1061ef376f51508c8f0e3;
mem[705] = 144'hfdd9f137f9670d4601c5f5d4fb06f63bfa21;
mem[706] = 144'hf1f50d78fd05fff80a30068bf87af4b10c61;
mem[707] = 144'hfa73fed40175f9cbf1a7fdcffb12f52b0857;
mem[708] = 144'hf608f41bf9870030fde5f45407470c900c4f;
mem[709] = 144'h0ca5fc19f0160edd05bdfbf901c5f2ca0168;
mem[710] = 144'h0064f34cf5d5f2f2058df00dfbfa0fd5f67c;
mem[711] = 144'hf03a065df940f6e3018a047e0c4ff6dafc16;
mem[712] = 144'hf6e0ff970028f18ffe53f367030cfda10024;
mem[713] = 144'h05ddf8fcf95af7680acdf331f81d00a8f251;
mem[714] = 144'hf51cf43cf4dd08e5014cf71efaf8083003ad;
mem[715] = 144'h08ff000f0e5b0901faeaf61ff70e0d8b081c;
mem[716] = 144'hf360fb5907b4f1ff06e2f3f5ff560140fe82;
mem[717] = 144'h074ff0af01d5f7400484f0f9f1a8fe800ad9;
mem[718] = 144'hfb25069df1f9014cffa6fdbd02d30e8dfee0;
mem[719] = 144'h0930064000f3f4bff2ec05c0014c00a607ee;
mem[720] = 144'h02d30654f9b20e9a0e70f701f8e2f9e50374;
mem[721] = 144'hfdb7f54902bbfaba04ad04d909b30aad023b;
mem[722] = 144'h04e4f9edf74f0fcef588017ff36a006bfd81;
mem[723] = 144'h012602eb0d29005d044afad4f47606f10231;
mem[724] = 144'hfee409b7061508d1007609f0ff95fec5f3d9;
mem[725] = 144'h03eef7980147038df9e9fb800185f403f478;
mem[726] = 144'h0751ff69f79b0905f407f4b2fed302b20c6d;
mem[727] = 144'h018303e90862ff06042c09e709ceff74fda9;
mem[728] = 144'h0870f043042602e2f0740d7afb92f528f5b3;
mem[729] = 144'hff4ef2fb058e0313073002ff0082fac90ec7;
mem[730] = 144'hf1a7094700070cff0b9efe1b0fdbfae5fddd;
mem[731] = 144'h0f47009ef2aafb5e0250fe0cfd1308ddf51f;
mem[732] = 144'h09220a340043f546fa9609d1f79d0d910bdb;
mem[733] = 144'hf3780c580c9bfbfe087b08c4015a0060f927;
mem[734] = 144'h0184fd330e01f3a40fe20b15f63affbef2c0;
mem[735] = 144'hf3c203ee0d72fa4d0e000743fa0fffd7faa7;
mem[736] = 144'h06b90825fb36030607180d9b028e01400ce6;
mem[737] = 144'h05a6f9f9f9780180f4c0f382fadc037cfffb;
mem[738] = 144'hf79cf2560120fd9e0b850bb2f1ddfd350c74;
mem[739] = 144'h0acb0f650d5cfc860c6dfe74f6e3f27103a3;
mem[740] = 144'hf57ff26e0417f94501ed0b0c0038035d0106;
mem[741] = 144'hfd62081d041f0993f932f5240eefff69fe33;
mem[742] = 144'hf8f8fbff0d5df880039df90007f5f68703c4;
mem[743] = 144'hfbab0ef0f452094df2af0d43f45af8e30cb9;
mem[744] = 144'h0c94f011fb12ffd5f7cb090503b6f6eff0ad;
mem[745] = 144'hf376fe1ff771061d025001d5034f027df921;
mem[746] = 144'hf85af4f4f5940cf2f54107b2007efc9d0153;
mem[747] = 144'hf6cc0fb4021006bdf6ecf96e0d8cf8dbfb0b;
mem[748] = 144'h0b7ff46cf46705280793f21efbb601dbfb08;
mem[749] = 144'h0d7e0c7e00060b56f35cfee8f8f6fb4ef83f;
mem[750] = 144'h098bf05d03d605b4fc7f02a508fbf8f50fc2;
mem[751] = 144'h09adf2a60c1cf5e6ff3a0d770fd50c5e090d;
mem[752] = 144'h0b0008b4fa5ffb47f40cfbf10f96f9520d34;
mem[753] = 144'h064409a9095202520a26024c0cc8f46ef0a8;
mem[754] = 144'h084008fcf9f8f88e0da207a403e50300f72c;
mem[755] = 144'hf7c60b1a03cb0fd8fb2008a301c9fc9a02d8;
mem[756] = 144'h00acf3f008d8019df7dbf34b0d70fa10f573;
mem[757] = 144'hf02e0ee1fc940e0afc46026ef3c40d85f489;
mem[758] = 144'h0f840119f29cf41d0601f43df82d0887f124;
mem[759] = 144'h0e4cf2850b4302c1057709a3fd18ff5cfa20;
mem[760] = 144'hffa6ff95f7e00e0604f50530fcecf0de0f1e;
mem[761] = 144'h047b072005d7f108f064f046f5acfaed0a60;
mem[762] = 144'hf1b2f118fcd9fc17fdf6f6da08f40b7a0d1e;
mem[763] = 144'hf3dd0bd7f9d30957068e01da0140f158f83c;
mem[764] = 144'hffd1f496f3930adef5daf1300c1f0ee7f7d4;
mem[765] = 144'hf3210ac2fc90f524f81df51d015bf0d2fbfa;
mem[766] = 144'h06f501d9f3f8f3f50669030e0b11fdf20d1f;
mem[767] = 144'hf5660724febafe2e0d000763f3d0097bf43a;
mem[768] = 144'hf8d8f3350e65f3a9ff250b80f0abff5e0dc2;
mem[769] = 144'h0036f87cf2500043ff2f09ff0918fe990ef1;
mem[770] = 144'hf991f42f06adff22f61df34d065ef8dd0980;
mem[771] = 144'hf09f0f410d22fe110555082ef1a30a1b03bb;
mem[772] = 144'h059b0bdf0bc60263f41b0830f6e5f4500ee6;
mem[773] = 144'h0efff3050228f27ff9d3061b044ef4500c05;
mem[774] = 144'h028a086206440e5f0854f14f05cf0fce0b2e;
mem[775] = 144'h07c4f63f093a0d3bf0fcfc17f59805e406b6;
mem[776] = 144'hfb7e099b0e70f02b0014f2c704c1010af214;
mem[777] = 144'hff16fc6b074bfa5709a90092f22f0a9d0b88;
mem[778] = 144'h0959f8280df5081cf6940398f0e8f34bf25e;
mem[779] = 144'hf51af428f386fd4df8a0f2e3f3ef0ba2ff6b;
mem[780] = 144'h0af7095b0c1f06c4f83909770b40f76cf2a2;
mem[781] = 144'h0db8fea9025b00c1f873077109760d050ad7;
mem[782] = 144'hfd640ad5f848f61afb6c0584f8e9083bf132;
mem[783] = 144'hf6bd0379fcdd003dfa120021f36cf8a0002b;
mem[784] = 144'h041f0607f1dc0e9e02a9f108f096fec0f94b;
mem[785] = 144'h0ab4f0b3f483f951f1b10358f6a509d4fdbc;
mem[786] = 144'hfd66fec402c9f525f19c0f15f8cc02f80b77;
mem[787] = 144'h0370fb090c9af4d8fe8a0fc1fd5a00f5f7ac;
mem[788] = 144'h0bcd05eff0d8f6860389fa47f4580db30e3e;
mem[789] = 144'h00f008f4f2a50e68fd260361f4b6f49e019a;
mem[790] = 144'h0dfe0244f6090a32f73f0cdef14cfa63f47a;
mem[791] = 144'hf3aa081205d1081001ca09ce0087f656098b;
mem[792] = 144'hf7150697f5490ed1fd360a3401f306ec05ee;
mem[793] = 144'h0ffa093bf2d703110ea6f86c0e640b910112;
mem[794] = 144'hf6170846f94cfe400663fa9df7c3fd53f5b7;
mem[795] = 144'hfbcdf73cf029f0210eaaff3501540e2d0499;
mem[796] = 144'hf6550a22082d0338f3caf02ff30dfa420875;
mem[797] = 144'hff180df1f3c6078f0148f179ffa2f380f04f;
mem[798] = 144'h05fdf3100280fd470fde0c0f0022f3acf590;
mem[799] = 144'h04cf025effa6f7ae08bff47f08e10e53fb84;
mem[800] = 144'h009708aefe0af0370151f8eef4cbf9feffc2;
mem[801] = 144'hf5aff57a03fdf82bf2f80b64f279fe3ff468;
mem[802] = 144'hf18ffdeef7a2f4f301510768fd460293fd9d;
mem[803] = 144'h0127f8d2fb0a08bffe17f65306b80e3f093f;
mem[804] = 144'h0838006103ad01b0037af799fe240ea7ffba;
mem[805] = 144'hfaadf5d5ffd8f7abfe330e0ef6a0fa6f0279;
mem[806] = 144'hf770f4fc09f9f3d3f6f20ea8fe4c077df741;
mem[807] = 144'hfa2700dafc6d09ba0f79f105f09af4e10f04;
mem[808] = 144'hf715f75f00df0a6408400fa0f607efe40d38;
mem[809] = 144'hfaca0459025d01aa08a3febf0589f83004d6;
mem[810] = 144'hfcbb0d2cf47d0609f7daf34406a5090c08a3;
mem[811] = 144'h0634fef1f2a20b7e068bf28b0c56f22900ab;
mem[812] = 144'hfcef0b44f8250e20fcd1f17ef6e9f109fb1f;
mem[813] = 144'hf6fbf053f1510b06fbe00e9ffa10f6790026;
mem[814] = 144'hfe7cf28f0f8d0967f76ef1e1f240016604b9;
mem[815] = 144'hf5ee08c2f0c0086d0ae607d3f9fe05700938;
mem[816] = 144'h0cde02ccf33104a7f221fbd4fcda06b1ffae;
mem[817] = 144'hf894f1eb0085fe20f7dcf4e3fdb7fb05f2a3;
mem[818] = 144'hf0fc035cf20cf896f04df071fbb4f3e402d7;
mem[819] = 144'hf73efa200fe207b7f08bfc030c23fa220694;
mem[820] = 144'h0f7e03baf658f6daf7840adef71b0fa8f55a;
mem[821] = 144'h02f0f04df2c1f6f3f766083cf11afe8f00fc;
mem[822] = 144'h0b09f649fa610765f07bfd930981080afc04;
mem[823] = 144'h03990cde0bc00743f87df68d090b0c000105;
mem[824] = 144'hf803fcf70fe70828f808f536f2a3fc0a0773;
mem[825] = 144'hf75cf0dcf71af84efab9f704075bf1270ec8;
mem[826] = 144'hf322f9970d3907e3f2b20a26fdf400aa0458;
mem[827] = 144'h0c82f3eb07e70f6ff01afed2fd1ef9100dcc;
mem[828] = 144'h01830558f7ff080f033406a107d5f25bf80d;
mem[829] = 144'h0f9af1ebff88fa26f2d802fefbbcfbe3084f;
mem[830] = 144'h02fe086c0c700d12f304f6ac01a70e16f1c7;
mem[831] = 144'h099ffad5f0100e2d0cb2f2c30eae09cb059a;
mem[832] = 144'hf169fd7b040af61e02fbfb46f06c0471fa3d;
mem[833] = 144'h043108a7fa1c0c1bf53b079807ce0a5705af;
mem[834] = 144'hf5f7f40cf019083a0a7d05bbf29df283f2ed;
mem[835] = 144'h0d6ffac40c7df2cd0b9006ad033f027f079c;
mem[836] = 144'hf7080aa40bac01920b71fd7cf78df72006bf;
mem[837] = 144'h0c7cfd1bf7f9f3800d5bf68008baf03a0b74;
mem[838] = 144'hfe75f0f7099cf7a602a7f4ed02160785f67f;
mem[839] = 144'hff53ff74f5ca0b0dfa7905c3046104b3fcd1;
mem[840] = 144'h008606790d18080ef7fc0d2d0744f7210adb;
mem[841] = 144'hf222f2a0f2c4f7cf07a30cb2022dfbc4fb6b;
mem[842] = 144'h0980f0a50d85f4d5f2f8f23affb3f4def48c;
mem[843] = 144'h0b6df67df184fe7afb8e020dfb9af1c8f872;
mem[844] = 144'hff720a2d0b7af9380b7dfeaefe03f4df0a72;
mem[845] = 144'hf639fffb03c601970675030300ff0625fc38;
mem[846] = 144'hf8e603760840fc7b0874fea90b9502450499;
mem[847] = 144'hfffdf024fdaffcb5f678f066f7ac0bdc07b8;
mem[848] = 144'h0dec0f57f494075d024ff3b2f00b085606a5;
mem[849] = 144'hfcda0ef208150f08fde006f4f57409b00582;
mem[850] = 144'hf8930317f5fb03690cfcff68f22ef0edf7dd;
mem[851] = 144'h0de00189fb99ff010e01f534fed2f616f468;
mem[852] = 144'hf589f0560db3f23bf3b0051ef8d0fbc60837;
mem[853] = 144'hfe5ff44df55901290a0d0363f806fcd70012;
mem[854] = 144'hf1caff900a1cf35f073f0f7c0339057f055b;
mem[855] = 144'hf59a0f17f6cd03860fbd03ad00c702470adb;
mem[856] = 144'hf58af94504dbf5a1ff9e034b00860d7f09a1;
mem[857] = 144'hf0ce0212f61cfa900f9ff655ffbcfede0a02;
mem[858] = 144'hfb1605bcf58905430f7003e0f5c4f4fc03ef;
mem[859] = 144'hf9cdfef2f5d40a64f267fb59f420f672038b;
mem[860] = 144'h0b280899f03bff95f1db06380b7a0497f9ad;
mem[861] = 144'hf7360c740b6df509fbbff1f0fd42fea6f870;
mem[862] = 144'h0beef096f283f1180b4cf63bf258ff0bfb8f;
mem[863] = 144'h0d760ca304d90500039df49e0232f39909d9;
mem[864] = 144'hf981077df6fdfd1e07ec04fdf9e90c20f255;
mem[865] = 144'h059bfc6b03a4f189f0340112081ff5ebf636;
mem[866] = 144'hf21ef43affb70ef10691f11cf3def5600300;
mem[867] = 144'hffa2f920090df95eff52fa5d0a17fc8df02c;
mem[868] = 144'h0d8600b40b1c0b880c3df125f46b06d2ff5b;
mem[869] = 144'h064b010cf10bf81c0e7306a00924f5c9078f;
mem[870] = 144'hf267f3befa25f7620baa0658080f0fb0f402;
mem[871] = 144'hf6bef73e0ecc03a1052d0b9df4420263f551;
mem[872] = 144'h04db0c39f434f9dc0f57f71f0088fbaaf365;
mem[873] = 144'hf53a0da50fd80c42f63c0521fc5efa9e05b6;
mem[874] = 144'h0d0a0f37f136f48e0f7108dff7c3fa31f2fe;
mem[875] = 144'h0655080efabafd86f89b04280cc9ff35073b;
mem[876] = 144'h0227f7e7f978f9fc07d3f374f300fa90f8e4;
mem[877] = 144'h0689f4fb0322fa780378fcd4f309f7700ce8;
mem[878] = 144'h0b6efbdbf70f0c71fc97051807c4fb75fcdb;
mem[879] = 144'hf4810d30f3eafa1d07d4fb64f0010c480cb6;
mem[880] = 144'hfefcf0a00ce0f8e9f2a20424f7a20ce3f0f4;
mem[881] = 144'h0d4d0a770487024af339fa14fc70feaf05b6;
mem[882] = 144'hfa72f37e03b808a7f7b2f3800596008c0077;
mem[883] = 144'h06480d37fa66fce3022a09cafa2d0ff5078a;
mem[884] = 144'h0cc4fc48f13df6a2fc7007b4f5a4f0ef0ac4;
mem[885] = 144'h0d13019f0bdb0aaf0a5f0b20034c0bb80b38;
mem[886] = 144'h090501a2f67309f8f24d05af0557fddf0ac2;
mem[887] = 144'hf57a06bafddff021f6cdfe6af886fbdfff16;
mem[888] = 144'hf4a4f1d0072d0dd8071905f0f0960c0406cc;
mem[889] = 144'hf6e5f48df019fe91f5bff6cbf22e0629f79b;
mem[890] = 144'hf609f7e3fc29056a0c21f042f200fac508a3;
mem[891] = 144'h0a0a0603f4aeff13f957fcf7f27a009ef670;
mem[892] = 144'h0b05ff2d0252f41e01720b9e090ff202081f;
mem[893] = 144'h015ff71a00c60373fa3908ebfacff57b0e6c;
mem[894] = 144'h0304f123f96c0a2bf658fc580c8cfe61ff10;
mem[895] = 144'hf5b9fd530c99f221080ef9be0a8b08effbfc;
mem[896] = 144'hf369f7f50b61f4fdfb1f01cafb4afbf6fc5d;
mem[897] = 144'hfe1b04c906a1f7100a03096cf1930846fd5c;
mem[898] = 144'hf161fdf0f3cf025002d4f25bf6eb0abb0d09;
mem[899] = 144'h006b056af4e8fdbf0fbaf6e5fbf0fafb09e9;
mem[900] = 144'hfc12f1e100def79bf9960fecfbea03150ac9;
mem[901] = 144'hf36205f1f19ef325f783ffa9f0be0155f396;
mem[902] = 144'hf334fbb1f529f633fdbafc76072e0673067a;
mem[903] = 144'h0f670367030901fb020b0cb10eb30835f54d;
mem[904] = 144'hfd2603b90440f8cdf4530657fea7f3230f3f;
mem[905] = 144'hfbbd0393fa18f181fe4204fefb84f95ef030;
mem[906] = 144'h017cfbc40835053a0848f7fe0d3bfcdd093d;
mem[907] = 144'h0368f2fcf116f63df9b204b108fdf693fca4;
mem[908] = 144'hfdc901120e450e62fefe0a0105bb0dcd0dd2;
mem[909] = 144'h008b0e7b07470d8d012e0b2df2a2fa0b09ed;
mem[910] = 144'hfa2cf5e302080683f79301ef0bec085f008f;
mem[911] = 144'h0dd009d20519f077002f057bf60804ea0a4c;
mem[912] = 144'h003ffc05f56ffbdaf27b059107fb0edcfc22;
mem[913] = 144'h0739076e0b69f6aafc650261fe3dfb1b0e0e;
mem[914] = 144'hf301f86cf404fe5a0dee0334f758f99a04fa;
mem[915] = 144'hf8f1090f07770bd0fcb2fa57f4300ce601ef;
mem[916] = 144'hf45f06dbfb9dfc2107f8fc0f0f93fb1f0239;
mem[917] = 144'hf6bb0bb7fead095b032d0b4c0cb20b74fd9b;
mem[918] = 144'h0f73fd120d080be5098b0f75fb920b95f934;
mem[919] = 144'hfffe002307ea0b42fb10f3de003bf177f698;
mem[920] = 144'h083402c909490b6003a80e0cffb9f07af2ae;
mem[921] = 144'h0c32fb6a06290407f0dcf8980833f7bdf381;
mem[922] = 144'hf4ce07f9000af0a6f3a50ef9f8b1fc16f8ac;
mem[923] = 144'hf94ffbe7f973f8ecf38c03900b40f5910a15;
mem[924] = 144'hfa96fa1101f6083dff2804d1056bf99806a9;
mem[925] = 144'h04e1f866f1f503ed086afac50a63f83afd3b;
mem[926] = 144'hf557effd0c0a0f86f002010201710cd10eb0;
mem[927] = 144'hfe32ff4afe1809dd09c10bfcf609f4ed08ad;
mem[928] = 144'h0f1302380723f2830c13f8f50cd8f98df3c5;
mem[929] = 144'hf8fbfd40faa602abf33fffbaf01af287097b;
mem[930] = 144'hf2300e29fa04f92b0ca1f772f042f5faffdb;
mem[931] = 144'hf045f5a1042b069df6f0feb904e1062cf1c4;
mem[932] = 144'hf48d08e6f238f92bf87500ec0b7bfe3d090a;
mem[933] = 144'hff6df07d036201f2014505d3fbb5f1a9f91a;
mem[934] = 144'hfff4f9c1068f084b00490ce20c96f20807f0;
mem[935] = 144'h0fd005680620fe70f15bf65effb5fc32fe34;
mem[936] = 144'hf83d093207ecffac07aef127f7b9f0d60a89;
mem[937] = 144'hf4e30a1ef8260deefa4efdbbf5c707f400da;
mem[938] = 144'hf69efc44ffe9f9b90d0b05800f890080025e;
mem[939] = 144'h0617fddbf37bf7770e5b0cd6011a077d0390;
mem[940] = 144'hfc87fb100146f201f6bb037ffa400c1bf52c;
mem[941] = 144'hf861044cf0b00ff0fd3409420445032f0094;
mem[942] = 144'h086e0aeef8e308eefe24039407e000d6f445;
mem[943] = 144'hfabaf1e80201f76a0d3bff26f4be0de80297;
mem[944] = 144'h06f7f7c60db3f4aef4a3f43ff7e2096f01d8;
mem[945] = 144'h07f804990d2101100e7f005af745fcf20992;
mem[946] = 144'h0cb50050f29407d7032af45b0708f1d90414;
mem[947] = 144'hf923f4610304f0420b93fb23f096f0bafa38;
mem[948] = 144'hf03706eef7f007e500bb0917077cf4acff38;
mem[949] = 144'h092d059bfb2cefce08a6f396fd08000e0b8b;
mem[950] = 144'h077bfb9df3c30bc6fcb9f4a40edcf5b90a98;
mem[951] = 144'hf7170d31fe07fa970c9b0c19f8d4022fff6d;
mem[952] = 144'hf7ae02eff0def400fac9f36e0a8ef4dcf8b8;
mem[953] = 144'h022001f4f9d20412fa3b0f48005cfd61fe08;
mem[954] = 144'h04c8fb4a04dff3befdc6f96d0cc00d980d6a;
mem[955] = 144'h0561f7a70d66fcae08a20ec2fcae0129ffeb;
mem[956] = 144'hfa00032bfe89fdfe04f10facfd2ef9d9049c;
mem[957] = 144'hff4e042df57df2d1f8740c56ff900bfe0c2b;
mem[958] = 144'hf0a70ee9f3050e30f278f578f25ef9850902;
mem[959] = 144'hf6bffb57003305f3f66ef3f1f191f7b6ff40;
mem[960] = 144'hf1760c0bf8d90a130a7bf9c40084ffc206bd;
mem[961] = 144'hfcf4fa4403e50598f021ffc1fdc300b20443;
mem[962] = 144'hf9ebfe2efd12f2f9094e00e601df0e35f2bd;
mem[963] = 144'h054bf1c3f7adf0be0604f253f775ff600dd7;
mem[964] = 144'h09daf3d5f1e3fa31f755f53002dff5a708e2;
mem[965] = 144'hfdfb0f76fe3601070bfa0dda0d69f48df208;
mem[966] = 144'hfb39f94c047ef0ccfec2fdccf04df01df8ae;
mem[967] = 144'h0fb9f53903b3f2a8f7d6fa57fa2506130f18;
mem[968] = 144'h088c0b120012036ef9c604660dc00484f186;
mem[969] = 144'h03970f82f96706cc0239f30d0a000766f78a;
mem[970] = 144'h0eae0938f4f802c50a5f02320529f0ebfada;
mem[971] = 144'hf7e0033c092ef14905b9fdafffdcf1280150;
mem[972] = 144'hf63a0d1df94f0950036cf0b0f020090cfae8;
mem[973] = 144'hfe9eff63ff64f12ef6bc0b950fb8f46bf580;
mem[974] = 144'hf67bfcaaf87ff05e0d53fa73f8b50053fabf;
mem[975] = 144'hfd94f75df170f48d0c6600e3f8c904420600;
mem[976] = 144'h082004e5086dfee3f9f2f327fbca0079fcca;
mem[977] = 144'hf0b8f085051008cfff9df718099508910239;
mem[978] = 144'h02eef9dff8f1f36a0ac10dc501a9f7cff149;
mem[979] = 144'hf4f603c9f908f795f57a002a0f5205a90b49;
mem[980] = 144'h0a64fa5bf767f36ff1cd0cd8f7a402a70cab;
mem[981] = 144'hf56c0f7c0976f6cafbc5f038fe6cfdf20390;
mem[982] = 144'hf22f0bedf4c4f798fbc8fcd6015b0baf00ca;
mem[983] = 144'h0a13f772f5480ca2f11af6530da3022d04ae;
mem[984] = 144'h0079f510fc070728f73208ca0f82092a016a;
mem[985] = 144'hfcc804e1025ef122fd0c08a5ff4efed40932;
mem[986] = 144'h07f5083d06a003a1f2e1f81d035d014b0233;
mem[987] = 144'hf9040ce0f2e0f5ee00de0f30fc0bf42bffc0;
mem[988] = 144'hfdbef4a401550d2d0f6208fef02df220f960;
mem[989] = 144'hf75c0371f37cf0bafeec06170c47011606e9;
mem[990] = 144'hf7a9058bfc30f348fe0df0bd07730d54ff03;
mem[991] = 144'hf255f1d60f2409e50f16f53e0fd3f8670e75;
mem[992] = 144'h031f09d404950d45fe51fb2d0c89f5f00fcd;
mem[993] = 144'hf782f3470bcd0720f582fcbd07e5012dff48;
mem[994] = 144'hfbebfed8040d078201df0383078703c507dc;
mem[995] = 144'hf71602af097a031ef021f88b0e23fccf05f6;
mem[996] = 144'h0d470bb60ddf09b90a5ef9b2f7c1fd680e89;
mem[997] = 144'h0becfe5209ee02b50a1cf5190e8ffe45fb00;
mem[998] = 144'h0a1e045cf265fd0e01e20dca067201eef01e;
mem[999] = 144'hf52208fc04affe37f44ff84e09cbfd090ec0;
mem[1000] = 144'h0e010e5d0c90028ef59af13d04c1fb69096d;
mem[1001] = 144'hf461f63afd8efe8805380ee6fb0ef30d01b1;
mem[1002] = 144'h0f2ff20e0204092ef973f1a1020efff807ce;
mem[1003] = 144'h09d0008b0bc5f4ee091500900eb6f2460adf;
mem[1004] = 144'h0bef042ff4090b30f285051c029cfc76059b;
mem[1005] = 144'h04820def04e0f73003b2fc38f5210ec5fba3;
mem[1006] = 144'hfdc806d5f511f713fc020e05033308ca00e1;
mem[1007] = 144'h08e505b806b5f92b0047070af9d6fffd0d2b;
mem[1008] = 144'h078bfb500c97f59205d9ffa80b8f0a950b93;
mem[1009] = 144'hf1bf083d0c2101bc0d3cf8c3f53b0dd50db3;
mem[1010] = 144'h0e4708b9f6e9fb31efe905ea0a37f67bfa2b;
mem[1011] = 144'h0bfafc0002ae0d8df569021b0f44f4cef549;
mem[1012] = 144'hfb2a059a09d0f810f3b405bcf09bf9aff433;
mem[1013] = 144'hf0b2fae8f978feb0068003fcf63efa0af868;
mem[1014] = 144'hf7ba07f307d5fcf20179fc990db0f2a307c0;
mem[1015] = 144'h0932f873f7e10c61f7cc011a0a63f9000883;
mem[1016] = 144'hff240505f5ae051cf0d905b9f7adfe41011a;
mem[1017] = 144'h0b71f28000cdf93ffd87f385091c023a0f81;
mem[1018] = 144'h0356f91e0a7f06b4fab0f5ddf783fc5b09d5;
mem[1019] = 144'hfbfd0cde009df28d003c0223f83e0bdbfd76;
mem[1020] = 144'h02ee0bcd0eecf486035e0ca9f1280814fd5f;
mem[1021] = 144'hfa2804c80c36f6db001af73bf247f06c085f;
mem[1022] = 144'hf4700c9df670f67b05f305a9f71c08300b8e;
mem[1023] = 144'h04440553fbdbf1b308170b18ff9a09f809d6;
mem[1024] = 144'hf55ff6220add08e20b9dfa60fd36f01a0791;
mem[1025] = 144'hfc3c0071fb92055ff14e094b05bb0d4108c4;
mem[1026] = 144'h07aef56704d50266f7e8f77bfc96f7bbf202;
mem[1027] = 144'h0357f0b9f99bfa80f66df0e1f22001db05bf;
mem[1028] = 144'hfe9cf7a8f137fff80139feb10a1efe8f040b;
mem[1029] = 144'hfb790f4df7b305e90621f67e09360d960233;
mem[1030] = 144'hf1cd0a27f62cf787f5c30993f113fd910ef5;
mem[1031] = 144'hfc0c06f3004a00b0fbfbf2440db006db0cbd;
mem[1032] = 144'hfab30be4f37c0b89f3edfd88ffadfc30f67d;
mem[1033] = 144'h075ef3f50d3b0eaa0e0005f6f333fe40ff61;
mem[1034] = 144'h02b40af009310df2f80bfc6df9f0f03d0ce5;
mem[1035] = 144'hfba30ad2fc1ef8c3f6550865008f0aeb02c0;
mem[1036] = 144'h0959011af24607070889070ef318fbd80bfe;
mem[1037] = 144'h06a0f297f5effb26f8c1084d0450060b0418;
mem[1038] = 144'hfd58fa04f3a306c404d3f99f0ffb09c70828;
mem[1039] = 144'hfef8f04dffae088b0333014bf6820d5706ca;
mem[1040] = 144'h0e69fd2c09e8f175f8ea0e6105a1051ff7be;
mem[1041] = 144'hfe850a7e0f6afac30a58fb2ef617040f07b5;
mem[1042] = 144'h0c5af080f60ff98efdcff68ef45307980d7d;
mem[1043] = 144'h04adf4fef970fe2b0cd70376f62c0e5df279;
mem[1044] = 144'h04a6f0e90ef2f14303f8050606d0fcec07f2;
mem[1045] = 144'h0b9aff85fc6ff7d6f78d05c50a9b0709f432;
mem[1046] = 144'hf1a309e0efe20c030584efd60d1ef1850f14;
mem[1047] = 144'hfff2027f021afe7c0dfc064308520935f0c7;
mem[1048] = 144'h079cf3b2fcdeffea09c0088204430ca9f997;
mem[1049] = 144'h069b0f69f12efd5fff91041c0adc058dfc90;
mem[1050] = 144'h0930f0b7f0c9ff6a087b0d7cfde50f520c45;
mem[1051] = 144'hf6c4f84affcef284ff73f146fe49ffef0e42;
mem[1052] = 144'hf13e08230d7af6a3f913f254f41dfdcbfe59;
mem[1053] = 144'hfd45fed2f2e6007efbb8f822f70e025e0a7d;
mem[1054] = 144'hf666077cf02e08a7f877f9800f09098c083e;
mem[1055] = 144'hf65afaea0d63060107c4fe600270f530f968;
mem[1056] = 144'hf36a05a4fd99f840f754f0e8051b051200cd;
mem[1057] = 144'hf68001faf2420f2b0876f5060b8dfb7ef7ed;
mem[1058] = 144'h030806a9f2fe06d6fdbff12ff63df4f3f1b0;
mem[1059] = 144'hf22f0012f72df32c0692fd82fd8c0eab01f3;
mem[1060] = 144'h058df8710dc103f8effc05da08cb0c8df61b;
mem[1061] = 144'h0781fa0df53f0dfdf455018c089c0428f448;
mem[1062] = 144'h06aefc5ef0a5f2d90488009b0248f6710535;
mem[1063] = 144'hf5e20c960717f072f103046506ad0c140dcf;
mem[1064] = 144'h037c083905ccf949f4a7fb71f1ad0e1b030d;
mem[1065] = 144'hf7e40ecafdb8f153079dfa8d03f2f919096a;
mem[1066] = 144'hfc0f0801fe500163007ff68ffef40c990967;
mem[1067] = 144'hf9910df3f7b806e4f2f8f1b3f5210b7bfa4d;
mem[1068] = 144'h0bfaff5b059d0f37f05afd61047cf52707c1;
mem[1069] = 144'h0e75f8b5fdd10d890a3beffb0d6ef41b0979;
mem[1070] = 144'h08eef6fbf1faf3e60205f219083f012d0b84;
mem[1071] = 144'hf16c0e4000a1ff91f1d4008a0908ffc00953;
mem[1072] = 144'hf5eff4defdf80719013f07e7075e099706ee;
mem[1073] = 144'h011303c6f9fb0bd5f8c3f8a5f212fe07fa02;
mem[1074] = 144'h060f035c0d63fb890bff0539070a0a55f22c;
mem[1075] = 144'hf6fc0930002c06e2f43804a6012f0fadfeb0;
mem[1076] = 144'h0f3a07f4f178fc65f53cf7c1f976fd75fe33;
mem[1077] = 144'h04e7fc1807f005fcf96208ebfc400e2e0de4;
mem[1078] = 144'hfd9cf164fcde05450a0806bcf474f49efd6e;
mem[1079] = 144'h05710399fa99f88efc0a0543f04f055bf7b1;
mem[1080] = 144'h03d2ffca08030ff00f20f654f2baf70d05ab;
mem[1081] = 144'h0e620bedf38903d3f526045ffb3a07330f58;
mem[1082] = 144'h092104abf978ff06f8f8f1cc012007490edb;
mem[1083] = 144'h064af7da027bf556f476fd6600be0001f3fd;
mem[1084] = 144'hf66d018ffc0b0c99f3b20cf608470f06f03f;
mem[1085] = 144'hfd44024af700f5b90e85fa2101bf0de1fe48;
mem[1086] = 144'hfe3cfc7ff835012405490813f7fdfab30a35;
mem[1087] = 144'hfdd6f7ab04330cba0635f59d03e10fe9f75f;
mem[1088] = 144'h0b7a04a60b40f962fc230faefceafebf0a24;
mem[1089] = 144'hfba3035401970a830b0af3cd0f0bff44fb26;
mem[1090] = 144'h015400ccfcaff3f10ccd0ed006310307f22a;
mem[1091] = 144'hfde7f987f61703e9003806f30ebcf6aef11b;
mem[1092] = 144'hffa4ffc30245f914f125f6f1fc2ff4930f60;
mem[1093] = 144'h03ed02bf0ef90577fadb027704430452075e;
mem[1094] = 144'hffca0487f70a0191f8d90087f273053c05ea;
mem[1095] = 144'hfae2fe53f9a2fbe4fa9507980eb70e63091d;
mem[1096] = 144'h014ff33af02a03b3f11afda00f4df118f67b;
mem[1097] = 144'hf1c7fcdc0edd098efd09f99508f7f59e0641;
mem[1098] = 144'h00e6f321f5a700c9087df13d03470ed6f0cf;
mem[1099] = 144'h047e08e602c0018f0093049607d50a430e92;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule