`timescale 1ns/1ns

module wt_mem4 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h0a6ae04411bdf1b4fb9714ea1a6af8d2eea9;
mem[1] = 144'h0effe663e9041197ee0b12d0fe3d19eb0118;
mem[2] = 144'h0300ec17f795f2f60bf308060fa7ebba11eb;
mem[3] = 144'h014f07ebf78aeecb0b771f40ff40f93ce253;
mem[4] = 144'he3d0faacf2b3f9810a0efba601a70836e105;
mem[5] = 144'hfad9eb0c05ecf3dbfacffda4e9f3e5ea0c62;
mem[6] = 144'hef8010ede5d41ab2ec0404dbf137f2570bb0;
mem[7] = 144'hf5f9f044ef50e916e258fc1004ed0f9a0b7b;
mem[8] = 144'h01bdee8a04bafe9fffd91611134119a40f40;
mem[9] = 144'h1ede00b8e87716c7eb56e1f41212f9691be8;
mem[10] = 144'hf31610bbe52de2f7086311be0059e5c119ef;
mem[11] = 144'heea7e9b8f2d20916120bef3bff02e674023e;
mem[12] = 144'h1f3af965f9c0eae8e4bc1ee6f0800bc8f9bd;
mem[13] = 144'h09c51ae0fc1b1ba012d0f071ea6904e71018;
mem[14] = 144'h137502421f401f11e58ce444e1dc134d1c1b;
mem[15] = 144'heba61bffe66214fde6e3ff611098eb6aec3a;
mem[16] = 144'hfce316bae8a0ef74f1eb155e0dc00eb7e8df;
mem[17] = 144'hffd3e8631214094cfe2011c2f3c9f74a0b07;
mem[18] = 144'hf210f8de156b193fffd2071a14dd0c7504cc;
mem[19] = 144'heccf1dd90e56fd2707a8f637fb7d0c280094;
mem[20] = 144'heaf2fc33fcf81c111c4815be05ca09fa0212;
mem[21] = 144'h16c406f305ddf97e19f6f4fbf40119d11644;
mem[22] = 144'h0e98e779f23cf7ece3af061105361ead1d8a;
mem[23] = 144'h0dcb16abf07ff4341a71e595f2f408f01579;
mem[24] = 144'h01241d911bce1f8c0b6bfeb9168ef9d3ef0f;
mem[25] = 144'he1ace7baf6cded54e0711202fd570eabfbee;
mem[26] = 144'h132fffa3151fe447105cea0c1ce00f89fd46;
mem[27] = 144'h0f0a144b17e002850307f5eaf5201ce30262;
mem[28] = 144'h133515cd0487e6b7f6aa0cc5148efb7a0f68;
mem[29] = 144'h1d140c0e185b024c00d2f497e199e33cee56;
mem[30] = 144'h0554176c01d008d7e3a20c6109c31450ed93;
mem[31] = 144'h1b1619c20552e915002d0c79f5a907c5e1e1;
mem[32] = 144'h133ae7851b09ef1c013cfff7069515cff1d5;
mem[33] = 144'hf97cf5d615a5e5fb164debff0f2df802e8af;
mem[34] = 144'h057c0232108beb25f03218c50ea11aace465;
mem[35] = 144'he8e5094de0ebf927195207e51e80fe9aeeca;
mem[36] = 144'h0d24105808d0151f1d07f5cee228f5deedc5;
mem[37] = 144'hfdf10a38fc8a0200186ef1d5e368e6771ea7;
mem[38] = 144'h196b041de28ff68f17ade8f3e7a9f630e4d9;
mem[39] = 144'hfdf91c4a1eb6ffa11e69fcbff3c500d2fb3c;
mem[40] = 144'h1a0e04410bec08f91b91fdcfea4a1207f0b0;
mem[41] = 144'hf77f0078f8ca07711ec40c2a1f88ee52e444;
mem[42] = 144'h063cf0b908f7fb91e612e8740ec5fcddfcfb;
mem[43] = 144'he779068a0beee27e00e21c360638e05d17aa;
mem[44] = 144'h14bb1b2e1c82fcf30f6c00b1f8650f4912c1;
mem[45] = 144'h0f3eef31157f10d501c80a5ffaceee811485;
mem[46] = 144'hecfdfefd17ebf57af092e3a004a104eefbfd;
mem[47] = 144'he5f7e911fc271d02e9a20a4ce97de568148b;
mem[48] = 144'h172f11def89af2251d00ea5807351aaf12e6;
mem[49] = 144'he5b1042df9b8f7f21dca1f2cff88fefbf009;
mem[50] = 144'hea2be773e64113f118171a21fe9808ade22e;
mem[51] = 144'h0c71089b17461dca0493eaf403551b55eba5;
mem[52] = 144'he79c1883e4531b43fb271ae605ef06d3090f;
mem[53] = 144'hfbc5141ddfc304cae7bd1c750463f369110b;
mem[54] = 144'h15351898f1611b6ff8d2178eeae1f86d0f76;
mem[55] = 144'he2371f2d0dd5fe06fb1c0513e96d1cef0262;
mem[56] = 144'h1d6605cef2c4e5b21a5ce34b130de6740040;
mem[57] = 144'h04d4fc0f104715e4e98812ecfff8e1cff2cf;
mem[58] = 144'he00117d3f21de98e0675fbbdf181f48619b5;
mem[59] = 144'hffa4f2a2e409ea7b035cea38f4bae3f71c14;
mem[60] = 144'h022ce5eb00aafeae18400b5b12c9e0380434;
mem[61] = 144'hf9821c89184d1c57f614edcc1a3bf2a4e8ad;
mem[62] = 144'h1ef01343e823195d038509e7176efacf175d;
mem[63] = 144'h11f210291e6a0eaf15fbe7251117115df975;
mem[64] = 144'h1997e9c0021c033defdbf6c2fb5afca91191;
mem[65] = 144'heeb2f38a1ce3ef5f14d9f97b08d418871360;
mem[66] = 144'h1e17176600e6f269159506811243e882e2d1;
mem[67] = 144'h0825092bff0a0e040886f346f7f5e427e3f8;
mem[68] = 144'hfc9bff9e120b1e62183a071a003ce3d71b0f;
mem[69] = 144'hf454e1ea0eecf32cfe21f417f720ff07e185;
mem[70] = 144'h09e3f4c1f14612dbed1711adfc6b065f0352;
mem[71] = 144'he9b418d7e390131418e211db12e516a6fc1c;
mem[72] = 144'h0adf06a0e5f91bf7f657eb1de2c9e400eea7;
mem[73] = 144'hff73ea9de6f71bb90f5e0203e6d0f40712c5;
mem[74] = 144'h142bf1cb077ee5b4eeea1cbbe1acf336102f;
mem[75] = 144'he5c2f089087b1028059d02190d861d7a161c;
mem[76] = 144'hebf9ee97e248f013e6721e48eebd0147fc90;
mem[77] = 144'h0323e66800e1167a03291bc9053612450f4e;
mem[78] = 144'he076f3b6e12ee41dede01849e7b40fbefed3;
mem[79] = 144'h15551610fdf81533e6d9fa7711a9e02d055b;
mem[80] = 144'h0a4ffe430bce057c00ad039e0648e724139c;
mem[81] = 144'he7f903e1f287f900eb17e233edc2ee200ca4;
mem[82] = 144'he624fbddf8cd1b29110b06dffbbee2b3f1e4;
mem[83] = 144'hed2e124f00fb1121e965054ff09a0b640bff;
mem[84] = 144'h1db901feea961b040075ff5ffea31112f0b2;
mem[85] = 144'h0c12eea00a7cf168046e04e7e8fd0e1a156d;
mem[86] = 144'h10f2e5bce04df37e09e3e02cedea07adef22;
mem[87] = 144'hfb0c0c1ef2cff8cfe3391e19002ae1d6f773;
mem[88] = 144'h124fe3fdedcdf32b13ca004cfe6d0c00edaf;
mem[89] = 144'h1ff2e970fe67ea22e94617700529ef69f2db;
mem[90] = 144'he3f20c3fe8cee048f0b6e97ef746eee5041a;
mem[91] = 144'h19dae2d904e4f74517bdfc4915c7e1b319ff;
mem[92] = 144'h1cbe13efecef068dfd74ecea08efebf80cc0;
mem[93] = 144'h17f4f9da1b1ae2520a4cf5ee0d08ea48e905;
mem[94] = 144'h1c4c1826ec111f2af3101e89faadfa04e3dd;
mem[95] = 144'h0eeef360eb95e19504e60a20ea50eea1ef7f;
mem[96] = 144'h0e0113040420156d00c814281b0c19e9e08a;
mem[97] = 144'hfc9801b8f00108db01a1f82bead90709e0e5;
mem[98] = 144'h197aeb031ea2f31ae80afe02f643f9aeeae9;
mem[99] = 144'h1ebbff6f15b21b57042fe6e41527023f0e72;
mem[100] = 144'hfd97e211ffb2fce2e12bfc77057c0e65f0ef;
mem[101] = 144'h1819029712740a3806cfe7fae837f460e9bb;
mem[102] = 144'hf2b0f15af40fe0f6f1b606d5130009b5ef29;
mem[103] = 144'hf4c010d71f090509ff06f6f4ee970f13ed1b;
mem[104] = 144'hfa22f0b5e5a31a570cd4020a0cfe0ef613a6;
mem[105] = 144'hfa160da8162de78c00c0f3a0e39ae955ec7d;
mem[106] = 144'hed31e32a0ba31bd004b6f9a4e40309670a67;
mem[107] = 144'h0912fd4c0421e503eae906b800d5e02cf52b;
mem[108] = 144'he14dfce412510a2f0cd5f670ee75fcdaecd6;
mem[109] = 144'hed370da3e8f2f559eacbe083efab189e177c;
mem[110] = 144'h0145135ffc43fb231ea2e8e408acef13e321;
mem[111] = 144'heb90eceae644e01b10e1eedb1ec5e3b2e940;
mem[112] = 144'hf0d4e87b0782fd48070c1c44e77de49916b2;
mem[113] = 144'h034916af188a1ac91bf5106c1c8f14030cc6;
mem[114] = 144'he3bde046f2ac0253e5ee062ae38b06250b4c;
mem[115] = 144'hfc04f9d2fa711072f9cd1319e47e011c162c;
mem[116] = 144'hffbe1003f096ecea11cdf9651eb2104d11f1;
mem[117] = 144'he034f9770faa106fef3e0ad9e24e15841c1c;
mem[118] = 144'h146219540a4f0fd116f6f6d717afe8ecf37a;
mem[119] = 144'h039c0348f249f6bf13d717eb1535eef814d1;
mem[120] = 144'h0c730d0d1224f7aa1e7202500d48e75e1c22;
mem[121] = 144'h0f09172b0ec4f76313dce05c1902f7cdeb53;
mem[122] = 144'hf65bf4c0feda0ec01c00fa36e9def81ee94d;
mem[123] = 144'hf45ef35d092cf7c9ff011e9ae9850c460579;
mem[124] = 144'he8300d8b08f9e1fffa2506dbe708f19e1403;
mem[125] = 144'he86f0c8f197b0c4dfb4de3d21c7e141ee618;
mem[126] = 144'heb16135119fde1ddf2f6eb4c02c00b5bf8dc;
mem[127] = 144'he8bce5790deff62b0fbe15feebbcf1e0039f;
mem[128] = 144'hfd15129918571e14fb7fe187f93d0e80faa3;
mem[129] = 144'hfe6af7c2eefcf3f0f9d303e5129de559fd30;
mem[130] = 144'he7e509c605ecf55d0a430e4d14741ae119c9;
mem[131] = 144'h15741829f9bef54ae3781806f1fdf061037d;
mem[132] = 144'he161108907cbf809f701e9b9f658ece4f9b9;
mem[133] = 144'hfb7c1068202c1aa9057aebf9f9ba14861b89;
mem[134] = 144'he4fa0b66006ff254f920f9410e7ff007ee69;
mem[135] = 144'hebcfe45fe520fd61fc81ea1ee74912070405;
mem[136] = 144'hf1fb1cc905f002371b59fa9c05701b53f037;
mem[137] = 144'h1961fea307ed153df0aaec14f1940836ebf3;
mem[138] = 144'hed7fe1520f07148e1c1c06151b910fc307c3;
mem[139] = 144'h09caf8f6ffc90f16020fed27e305fa94e559;
mem[140] = 144'h09e90061e610e917ebce0317e57a1b14068c;
mem[141] = 144'h0df9e1ce19bae5f9ee3fe87cf174f8b703ed;
mem[142] = 144'hfd8104c31c2fe641e249e93dff870f1b0209;
mem[143] = 144'h09f6057a0e17ed05f5c5ec2105a313c4e32f;
mem[144] = 144'h1559187112cd174c1424129a12ac123aed17;
mem[145] = 144'hf2b01c2bfe6104b1045cf430fc79110712c3;
mem[146] = 144'h085ef7a90491ef30f82cfa1ee6c9f2cdf687;
mem[147] = 144'h02820d531cf9185be8b409730386169515ea;
mem[148] = 144'hec4e0559fd410f90164f17b1f0b4f4ba18bc;
mem[149] = 144'hf5b1153f114ffea5f792eb641e49f365e6d2;
mem[150] = 144'h1a2bffe318331b640e6af962e8430c37ea4d;
mem[151] = 144'hedc104ccf700f96702d2142a1ff50b681af6;
mem[152] = 144'he8c3f4d2f487075ce6030395f8bbe51415d3;
mem[153] = 144'hffc1ff3b1ffb1d22eb451a50fe451170122e;
mem[154] = 144'hedade703f80ae90be9f2fb17f577eb2602cc;
mem[155] = 144'h088af343e5b4167115770d2618130f280f94;
mem[156] = 144'h17bb0a37ed971ffa0b90e89204491da40419;
mem[157] = 144'hf223e4aa07fd1881093b0a16ff361578e21c;
mem[158] = 144'hf83a027a040df51af4c1f028fcf3e4d01426;
mem[159] = 144'h0eddf568e6a615a3fb71130002bb11b1e842;
mem[160] = 144'h014be5bc102e1b931fd1093f19fb0f470233;
mem[161] = 144'h052be0eff2b1f6bdebff0f68eb05eee5fc46;
mem[162] = 144'hf7b0f812076a02e5e6e6063fe06302e2e669;
mem[163] = 144'he19c14e5f57201a4f8fee386079d14afe321;
mem[164] = 144'h197bf7b0f05919acfbb7ff1505c20637fcf1;
mem[165] = 144'h124903d6184317b3f14213da18f7141117ef;
mem[166] = 144'h1fdafd7ce4dee05ff215fad7e60df86518fd;
mem[167] = 144'h042decc1f512e978fdeaf2771087ea651050;
mem[168] = 144'he0c3fa82081dfb5de8a70b3de2f0e5cce100;
mem[169] = 144'h04da0113176f1566f342194c0dd8fec40176;
mem[170] = 144'hf512edbeffba0ce5ea1e19d0f54213be1bae;
mem[171] = 144'heaf4e18301b3f2bb1a36fa66083ef63a1558;
mem[172] = 144'h1ce51a2601dfe833fe7c081917261315facb;
mem[173] = 144'h0c4005b6193ffe24e69bec0000ca16ca0dfe;
mem[174] = 144'h048f1262071f0aeff773eb4e06f614131ee9;
mem[175] = 144'h02080a51eb06effff27402bae212fc05fe76;
mem[176] = 144'h1599e4c7e3b3f1c6fe4ff922eb560d8deb54;
mem[177] = 144'h04cb05af0f37e80305e1fe34fe83e418f1f0;
mem[178] = 144'hf474fc3f03e6e6e407edfb3ff199120412bf;
mem[179] = 144'he070e0afe890f11cfd491c11fa3ae10f1090;
mem[180] = 144'hf8eaff7d0234171206c517090fb41e89ffcf;
mem[181] = 144'h115a041df603e5651f9ce3cf0661e16bf999;
mem[182] = 144'hface03251dd8fe83f91414eee5fc03cb1206;
mem[183] = 144'h1a2701210848ea46e7f6e3510126efdc139c;
mem[184] = 144'he2510b7e19cee865e3b600bd052b12d2e8bd;
mem[185] = 144'h0f20f6b9e3f5e55fe66e15c80329e33410ea;
mem[186] = 144'hf1941b430e530cbfef77e093febfe0fbdff3;
mem[187] = 144'h0ddce65df16e0a59e01c0f960988fa5a1811;
mem[188] = 144'h1d3ffe02068d002d17e1e5d9e8031498f348;
mem[189] = 144'hec5cf17f0da90e6f0f721da8f308ee69f320;
mem[190] = 144'he6ae008d1909194e0577ed1ff8bb023a10f9;
mem[191] = 144'hfcdae737f00d0d94000a1c50e1baf9981cc0;
mem[192] = 144'h0c73fd0d1fb01c1af324e28ae75a1fd50826;
mem[193] = 144'h1bb1026c0b271ee21459062b1a60e58a11e2;
mem[194] = 144'h12ed0108f1e9e8c707c8e7cc1c56f4f4fdfb;
mem[195] = 144'h124fe61e0c82eac4f53ee3b6f08afe610b43;
mem[196] = 144'he68801bde5dd1e4af82a0e9be53ffce4f7df;
mem[197] = 144'h0a24064b13cc0b1d09750554f96c1593e8df;
mem[198] = 144'hf105f52ae881e8d1f1e70e78ec7deca21849;
mem[199] = 144'h0ccb1ce4fa77e153f001ec0efe811e670770;
mem[200] = 144'hf695e077f09109cb07410428f1cee76b1625;
mem[201] = 144'h15a5ec99eb560714f63cf080ecff1873fb1b;
mem[202] = 144'h0ee20bfa1f35f7d413250b400ca10610e556;
mem[203] = 144'h0bae04e71cd71d62edb70ad90ab206d91b83;
mem[204] = 144'h031311a4e0f80577f26808e20eaeeefae819;
mem[205] = 144'h06afe7271e260ba6e742e55bfe4f08091e04;
mem[206] = 144'hf5ac1e8b00621877eae7f050e12bec9bfd05;
mem[207] = 144'h071aee051069eaa30c6807f21146efa403b9;
mem[208] = 144'hec9c00e4edbafc49e20efaf7e1f90cd9f3c8;
mem[209] = 144'h12bbeca3f3c3f81ffb4d0821f919f26ee699;
mem[210] = 144'hf34ff334e9b7e6091a58f6660b26e6130bfa;
mem[211] = 144'hfca202c51b0ee2e116dceff0faac1c6b17f5;
mem[212] = 144'hf661fcb803f0e9b20e2c02b9f7ffffc3f86e;
mem[213] = 144'hf90004361e2d0f55f8e30cf5e133ff39128d;
mem[214] = 144'hf0a3ebec0624f23b043019effc5112141335;
mem[215] = 144'h18abe78c04f9fdcafc810b3cf16c114b0b62;
mem[216] = 144'h136ffbc8f90a1136151be607f3ade031f406;
mem[217] = 144'h0966f4801031ecf002a9ed5bff7af7e41388;
mem[218] = 144'h0d46f76c15400465008b1c10f65ef3300981;
mem[219] = 144'heb87fa1de49305a8f098eb75e46cedcdf2cc;
mem[220] = 144'he751ec36f416e7b3066dffe3ec140503042b;
mem[221] = 144'h0890eaecf853e1fee6a2ef42e09e1ec215e4;
mem[222] = 144'hec910971edbc17e0e3e1fe01fd5bea40ef33;
mem[223] = 144'h0b02063ae8a9f04ee8a71350ee05ea8eff9c;
mem[224] = 144'he2f817bd1116e9920f81f6caf4650f331946;
mem[225] = 144'he607e376f53ee2c7ede9fe18f749eded10b7;
mem[226] = 144'h06e1fe9d0eeaf3e606cb02fef8affc450bb8;
mem[227] = 144'hf27b16ccff34eaee06dcf802f874fd5af52e;
mem[228] = 144'heb6de91d168ae7e2f43c085ee5921e30fd51;
mem[229] = 144'hef3bfe93ef2cf8a4e76a19dd116ce692e882;
mem[230] = 144'hf5c4e75ff83c0271f8211217f46307b6e557;
mem[231] = 144'h0f911dfefe9001f9ec100b211da416431f29;
mem[232] = 144'hfbe106cdec97018c060afe1600efe116033e;
mem[233] = 144'hfcb61239e06305a9e5b1f6490a83fb7d1bf3;
mem[234] = 144'hf25c1f921fc5f7c71e7508afefdbea42fd57;
mem[235] = 144'he635eec6ec4ee075094ffeecfc250b08e77c;
mem[236] = 144'h131df334f1ece186faf0f880eae401470ffe;
mem[237] = 144'h014f083012e3e06c1a15e73cfc82f98ae533;
mem[238] = 144'hef3708ad0cf3072ce8110d1beb91f6b715bd;
mem[239] = 144'hfc20f6c0e716e2c108791e6df1520120f7fc;
mem[240] = 144'h155ef2351efcfad1e2331f201702e6b5f78c;
mem[241] = 144'h1109e974e7c2e9ee1d03fcbfea9ae977f7df;
mem[242] = 144'hfd91e066e28a1402ff10e82216d8e1dcfaf9;
mem[243] = 144'h173ef0eb005d1b40ec9efa77e62a1666012f;
mem[244] = 144'heff109c70e8fec671cc2f139f45d10d50df0;
mem[245] = 144'he7d9f5d0fb0d0a1df3b2f2870c76050dff16;
mem[246] = 144'h1278057ff97bf59ae848f4ec093beeb3ea6f;
mem[247] = 144'hfc7617150cff02fe09600541f472f7a8e0ee;
mem[248] = 144'he93a18e61474078cf704eac1f5fb046d1379;
mem[249] = 144'hf2bfe3ec0fe71b3308edfb9ce77bed38ff3b;
mem[250] = 144'he06ae41e1e3a07a7e60c04bc16abe12bf670;
mem[251] = 144'hebe4f839127cf3b51d3616ecf6841a0eeffc;
mem[252] = 144'h1175f14d13131cc512130277ea9d14a0fc84;
mem[253] = 144'hf3acf0fff6faf3c9014d1e8be89f0ad20564;
mem[254] = 144'hf110174413a0fe780c38f02c0d681b440a52;
mem[255] = 144'hfe0dfc6c018d1bb30b48e7f0f0aceaaa179c;
mem[256] = 144'he60f0fa6e9dc1aeeea44f2fcf56a09c71698;
mem[257] = 144'h0a4ee0cf1413f720fc480ff504b704f90da2;
mem[258] = 144'hf2baeaf9134e00de04e9e5370b300b3a0a33;
mem[259] = 144'h0a0011a3e04ce6f4e92fea92e8670246fd0d;
mem[260] = 144'h09060b2e027af07d166205e0fd021eb40eb8;
mem[261] = 144'hed6713f21fbfe132e2981706e292e9931057;
mem[262] = 144'h08bdf75012711411e9c4ece80f6de5ace1ad;
mem[263] = 144'he797e39b1b0ce2b0eee8e87dfcf90b47eeba;
mem[264] = 144'hf3f705b0e3a1f4651e390e2612781d65e12a;
mem[265] = 144'he5bf06730d68f9d500e9063dee1e0d6cf752;
mem[266] = 144'hf3af00cd07030c7ff502009e187614bfffa5;
mem[267] = 144'h187f08efe60bfa8713d1fe02f09a1e3710f5;
mem[268] = 144'h1188fe80072d08670361f2f613340cd31961;
mem[269] = 144'hf5ceebd113d41c820429f1d31e7b11b9f812;
mem[270] = 144'hfe47e4920af4e258fb14f3fff32ffe8debce;
mem[271] = 144'h1cf31fe91368e69af7501bb2eab3e8f00be8;
mem[272] = 144'hfe721e05e9e1faa1e10ef478fe721aec0385;
mem[273] = 144'h1af40669fc8b1b28eaf50f90f61eeb7c1961;
mem[274] = 144'h1546f36dfa0117741edaf28606ebe7200888;
mem[275] = 144'hf23808d3ec0f1562111b1c490708fbc7eb7c;
mem[276] = 144'h1e730ffc0afc0e9a11a31772ea4fecfbf583;
mem[277] = 144'h07d2130306dd057af7b0fa280efc1b011d1c;
mem[278] = 144'h0fd2e4c1023901680d4509ecf54c1ea3f47a;
mem[279] = 144'h1c1d13cef35c13c8e8d80c36021efb7df508;
mem[280] = 144'he8191007fcde05d3f0d31edb110ce7c9f3f3;
mem[281] = 144'h0e0c1051f3df1c09e0abf827fc150236faab;
mem[282] = 144'hf5c41386efeff74e1f90f88917980decef50;
mem[283] = 144'hf133ea14f5a0f66c0714fab5e2f81fae0085;
mem[284] = 144'h0cf81f4dff780933e120e950fd9a051ff31d;
mem[285] = 144'he41bf8fd12621be6fe751820fb1f0497ed01;
mem[286] = 144'h1ea5ede901e2e8ec0e51f66de1671f0bff5b;
mem[287] = 144'h075de9de05f41b15078ae8a0e013fcd5f529;
mem[288] = 144'hea7916d4f3e80394f3f9031b1c6b0c030b9e;
mem[289] = 144'hf0f503841680f2c70531e633e3cbe017f762;
mem[290] = 144'h04830fa5151f1ec001300b51fc20ecc7019c;
mem[291] = 144'h09410e6711e6e9b709c6e83209ffe190163c;
mem[292] = 144'h1aecf3941715ee4cf32b1b3ce3d5e207fdb7;
mem[293] = 144'h05e9f20fe11bf5430e4f1fdf13ed0e801c30;
mem[294] = 144'h19cef526fcfcebe9f123e6f8144c0965ed1a;
mem[295] = 144'h062cf18e024d09d4e350e136122309d3efc5;
mem[296] = 144'h15befa5defcd17da1e401ad0f0a6e5fbfbff;
mem[297] = 144'h18c8114f1e3c0f590df01dc70c3411b8f8e6;
mem[298] = 144'hfc690ebc1d5df844ffa71797eb261144f372;
mem[299] = 144'h1baeedfd08521e0cf52e0abb184be8350c9f;
mem[300] = 144'h1191e3e6fa480cb9f53b09eb178dfe8f0667;
mem[301] = 144'h0ad91000e19d091f0f6111a9f947fdc5fdc7;
mem[302] = 144'he0561c451a70160909150823e7f9fbe0083d;
mem[303] = 144'h0c901f2eef06134c004fe08010aafa88ed31;
mem[304] = 144'hf4bd0ccce97de90f0b3ff416e227eabff200;
mem[305] = 144'hfcee062dfc070a8b097aff0de157e01a089c;
mem[306] = 144'he483052e1e2af4e8f652fd401d8601f0ec42;
mem[307] = 144'hf0df1942071816c7f5e9105815d30048e2f9;
mem[308] = 144'he372137a0353063617da1cdffc79ea1ff82c;
mem[309] = 144'h1ddced9c1d46e77f11c50769e425e8f5f415;
mem[310] = 144'h200005ebe0fa1855157218b4f02c0e5f0214;
mem[311] = 144'hf530e12d0b4605ed116fe727fa610b62fdf6;
mem[312] = 144'hfc8f179cf7e31ac7033dfa02f75409c2e076;
mem[313] = 144'h0916ef37062fe43b0c67f4c8fd06e93e0a62;
mem[314] = 144'hecbd063d1d28f689fda80751ee331e61e51b;
mem[315] = 144'hf312f2ebeb97165dfa58070df5c31f52f1c3;
mem[316] = 144'he03fe6b702a9f59f1037e12ef34af797eb68;
mem[317] = 144'h0c591b60ee8f03a2fcd6e53f04851661f2b8;
mem[318] = 144'h10090b92f369e16007dee3e3004be0d8e2e5;
mem[319] = 144'h0f6f02a2014b0e930bb9ed741f0ef326121b;
mem[320] = 144'he648ee95138611acf3ce0e41086f12c5faa2;
mem[321] = 144'h1fb6ee61f659f1f1f5271aa006fbffff053e;
mem[322] = 144'hf10b0ce0fb09ee0e1ee7fff314aa082200be;
mem[323] = 144'heb2f112612b7064ee39e08f8fffd18170182;
mem[324] = 144'h19ccf3331a49eb24f801e445f2420e10e418;
mem[325] = 144'h00f3f002e36c0a8de6681d6cff24ed491b18;
mem[326] = 144'h1e8a0019f44fe38beaeb059607460748e220;
mem[327] = 144'hf2c0f6aa141f0e170d3e1cd51a361c93eae5;
mem[328] = 144'he65009a4ea0ff2c6fc7b0fc6f154edd0fcc1;
mem[329] = 144'h01a10c7afcb6e93204e404fd1baef0ff1df4;
mem[330] = 144'hf7a5e7350a591129fd3d0cdefbf6f3bc1999;
mem[331] = 144'h12980bb40d51f42905681fa7ed2d12b1e42e;
mem[332] = 144'h13faf46ae73d0fb40b610795f0fe180ce2c8;
mem[333] = 144'hf9451bcf1e100a6d16db00f1e577f6c605a4;
mem[334] = 144'h19fdf52df38ded56e8c310421c92f5560436;
mem[335] = 144'hfc51e11b01bcf65bfb6518e400ed0052199e;
mem[336] = 144'h1f5ce2df01171c6d088ff29a1406114503c7;
mem[337] = 144'hee5614c6e4c3e7660c6505e31fd4f2250b2f;
mem[338] = 144'heaf01380e373012b1f7de3bee0acf7e90fe4;
mem[339] = 144'hf797ed3d15a0eca8fae7f3a0f3a91a21eee5;
mem[340] = 144'hec29f18b03a204d013191c8eecbf11bf1ee5;
mem[341] = 144'h1c3beda91dfb02bd1ae0e27b1f96ff7e0819;
mem[342] = 144'hfe761201f17902660b56120116d21e7cea15;
mem[343] = 144'h0043087c0d85f968078bf05be7b900691c94;
mem[344] = 144'h1c4f054805b005ac1980fc18ff6cefaf03a0;
mem[345] = 144'hec0af4f81393177413b8e99a1178011a100d;
mem[346] = 144'h0fd402fbfa2be7071eff1d1fe2f5f1940453;
mem[347] = 144'hee9b142cfe76f7a2f6a1f79ce54d06701bd2;
mem[348] = 144'he339108401120986fd06e894ee58ebf0e14a;
mem[349] = 144'h00d8fd600a7d1a98f75a0648f0affc24fef9;
mem[350] = 144'he4abfb4c014109e7f67201eb109bf16ae830;
mem[351] = 144'hfc9c1489f09d16b601c30cb90465e07a1dcb;
mem[352] = 144'h1936f572f6c912bcef8be5810092f65b1561;
mem[353] = 144'hfea5f2a7eac716d5fbae0783ea9c01540d54;
mem[354] = 144'h03dc1687125ff698195be4b6e91006d0fade;
mem[355] = 144'h0267e2c60bfe130bfd7fe768eaddf24119cf;
mem[356] = 144'h1f87f15016effd601446ffc900a10947062a;
mem[357] = 144'heec8036dfa8deb700bfeeb8df8f1f2a90920;
mem[358] = 144'hfe9314aff9b9086fef8e062feb76f00806e9;
mem[359] = 144'h1611f72a1197edc202d01d0417d6fc5cf736;
mem[360] = 144'h1d9ce2850395fa7e0027164dfd1ceb96efa3;
mem[361] = 144'hf0581b55fb7ff4a3e26c08dfe0a7f91c05e7;
mem[362] = 144'hf46b18d8e6050ac3f5b3ee9d08191891e855;
mem[363] = 144'h1501f2f91357ec4ef97e16c9fc3cff45e9f2;
mem[364] = 144'h1c3509cee9411c6fe33d1e661c2ffbd8f1da;
mem[365] = 144'hff1ef46aee9de448e37c00d4e0c8fd4419ae;
mem[366] = 144'h0a4404cff850ea5e1a0a0efa06b7fb6de252;
mem[367] = 144'hee3be353123803b9f858101be58ef2b316b9;
mem[368] = 144'hf7ef1a25f158fe86fe2d144f1e22f726e4a4;
mem[369] = 144'hf247e44e09d8f07602c5013e0acb1bdefa67;
mem[370] = 144'hecefe789085317020f76f5a0fee6162b0f33;
mem[371] = 144'h1b4ae9d4e536126502461d28e31fe87e02a4;
mem[372] = 144'hf4e510ddfcfa18821ff0e45be13ff5a3fccf;
mem[373] = 144'h03c901a8168bf964e739e70b0cea0a830745;
mem[374] = 144'he464196ceeb71858096deb2b0048f1fb0512;
mem[375] = 144'h1c8600d816ff081ce210007a09b0e633e592;
mem[376] = 144'hf19b0823e93504611acffc821a9219af0544;
mem[377] = 144'h032e0078edfd10d3f48207181b4ce85f1e9e;
mem[378] = 144'h1e9cf055e6b11a0d0b8c0e92e5e2fa7cffe9;
mem[379] = 144'h1e3eea50e69d0623e02812f9fa0d0c710b7e;
mem[380] = 144'he9e5fa1af97de114132de6681690fb41f7d4;
mem[381] = 144'he1a2e716e82af97f1bc91add0bcf017cf0d5;
mem[382] = 144'hfa54fd57fac71410e4a9fdd20c960c71fbeb;
mem[383] = 144'h0c5411a40cc815eae34cedccf404e271ee08;
mem[384] = 144'he1e10db205fd045d07fd0ebf1791f8fd1ddf;
mem[385] = 144'h099df0ea1c92eab307ebf8cb1648f2de0e39;
mem[386] = 144'hff830a110095f0a40a8bf58205290cf10bfc;
mem[387] = 144'h0ff20df91398e61f150614bfee74e003e652;
mem[388] = 144'hee90f464ea48e06be2e3e9d5152009e61e35;
mem[389] = 144'he560f38918c9ff6d1023eba6edc6e69fe322;
mem[390] = 144'hf38104650bbd1031f564e5260d8c032e02ef;
mem[391] = 144'h164b1fecf1ae14510495fc0efba4fcaf1e32;
mem[392] = 144'h160af99f1ec210d81bb40dd61293fbc1082c;
mem[393] = 144'hf4eeefbdf6bb185cfa8cf5c2e698e6fb0365;
mem[394] = 144'h1d6df9511d931318f7c3ecbd04ddfe8eff1c;
mem[395] = 144'hef1014f308e1fed60b3debe11f53e3b3025e;
mem[396] = 144'h0e8ee845f46af9fa130c1686047b14fc196f;
mem[397] = 144'hf447e33a0ef2eaad0061e1e40cc906700be4;
mem[398] = 144'he065e1fc0d3e1242f2031fe71d450d7a061c;
mem[399] = 144'h1539f440fcc415c21fa314620b7407d90a2a;
mem[400] = 144'hf51c1e040624189d0d0df36aef4914d5ec65;
mem[401] = 144'h1a79193a1c670115fdfee357fdc8e78c1736;
mem[402] = 144'h0eae1030045515ff0eef1f0af2bff9211d27;
mem[403] = 144'he974e83be8a0eaf91fe5e9bcf77cf45916da;
mem[404] = 144'h1c66f6d9ef2ff784ef28f2f3ecd3e2ec0c13;
mem[405] = 144'h14c5155afee2fc1a0fda187effed10fc0ab1;
mem[406] = 144'h1b14e28bf752f7e3fda5150aeebc1d0a1d46;
mem[407] = 144'h02d10dfaeba6046d1d67efc7e8bd1431f061;
mem[408] = 144'h1844edb20f200613e7580a0a0863fd15f7a9;
mem[409] = 144'hea5be687061f00561710e1a8fa2fe78e1070;
mem[410] = 144'h163ff04b1b51ed41125efc410a1b0e9efb3c;
mem[411] = 144'h1d1cfe1ee400eb451b19f6ece9580acf1d83;
mem[412] = 144'he9e61748f25c1bb60f4c0a3be23409faeaba;
mem[413] = 144'hf6c8184309ac07381bd0e78ff40913781cd8;
mem[414] = 144'h06cce88cfe0bf83b1dd61bd31c5fe2d51765;
mem[415] = 144'h049b0b5e0447f78b07f5192301c0e499eacd;
mem[416] = 144'hf97ee128eba607921a531bedf60705b01da0;
mem[417] = 144'h14f4f5f0055df085055ef2f1eb6b1129ffc2;
mem[418] = 144'h1d1f0cf0f3ca054dfbe6101bfc160499f3b5;
mem[419] = 144'he02fee2104790694f879f925045801ede2bc;
mem[420] = 144'h13e50b3b0727ea6afb94eacdfb4d1785ff3b;
mem[421] = 144'heb3ae518e5c708aa1456075fe38ff2db1dd2;
mem[422] = 144'h0bea1d47ec5516330d38e9d213b4f01e0861;
mem[423] = 144'h015517fef65b0d16151a1785e12efa6de324;
mem[424] = 144'h0800fda5e6d9fa3a0f38e44ffef0ec15e610;
mem[425] = 144'h1a5b11b60866fe2109280ec7e4501c9af140;
mem[426] = 144'h05affafe16660415e35af5b2013be9a9f96f;
mem[427] = 144'hebc110d21303e2ea1f89e66815c61f80f8e6;
mem[428] = 144'he40fe5e0f5831af011f9e9070126f70c0b44;
mem[429] = 144'h1bb502d4f5ca19cbf653e9680973e1b8f3bf;
mem[430] = 144'hedea00631c15e4ef01e20098f230e9050150;
mem[431] = 144'h1963e52eea790bf7f637e050e9d0e9de0088;
mem[432] = 144'h17bef52614821143f79d070ae2fae94e1e32;
mem[433] = 144'h1fd9e95af8440adbe68f06fcfd280653e2bc;
mem[434] = 144'h10cb06ba0fd10e0bf9940961f97deffcf5e8;
mem[435] = 144'he821fd0704c8f4ceec2afd9e04761511e917;
mem[436] = 144'h1b2ae225fbc2e4e216390f0d0eebe697f6df;
mem[437] = 144'h0411f9a7ff48e9850656107fe245ea4e1b02;
mem[438] = 144'hf254198ee7a4ff96f6d3e3ef050d0272065c;
mem[439] = 144'h01adfb4a1b270e49f917f8ebf768065fe609;
mem[440] = 144'hfd8b0befe5d01a640a5b0745f3551b890f5a;
mem[441] = 144'h1589196bee9b0bd5f948f76e0e80f4f21657;
mem[442] = 144'he6ff0ae8e0f00659e7180ad1e479fab8fc90;
mem[443] = 144'h0f521893f64df8d1eef61c11f495f4e91617;
mem[444] = 144'hf8a20e691d740f53e53616831ec7f9cd1208;
mem[445] = 144'hf17c0635ecda0c180b2109d904c2f9def3e0;
mem[446] = 144'hebedffe0108c0df407910081edd70eb21fec;
mem[447] = 144'hf5bf00dafaa5193b12f3e7a7fda7e856f23f;
mem[448] = 144'h006d0085f21be760e91b0a620456e53f1106;
mem[449] = 144'h0dae088200ece99bfccf1e2ff729ff6f0bf8;
mem[450] = 144'he520e273f58cf5fcedf21881e8ca0e8df8c5;
mem[451] = 144'h1aaffdc7e108f11b1f830f3811d70b1cedeb;
mem[452] = 144'h0dfce99a06dc19acf8bb184d01b71c9bfb9d;
mem[453] = 144'h1410199a08241b18044702dfff51f069fa98;
mem[454] = 144'hfbc5e9c009b0e871f3af05c11e9f054de30f;
mem[455] = 144'h0801fdbcf85408e613eee5cfe11ce58cfc3b;
mem[456] = 144'h0c56f14601bfea711103ef1d198e12e20ce1;
mem[457] = 144'h0b13015de12ef2e0f84ffbb61c75e2680707;
mem[458] = 144'hec601b14ff0a029f0fce1edf1809ef021039;
mem[459] = 144'hed52063e0d62e16017eee48f0097e50ce631;
mem[460] = 144'hfd4be4ff0325ec2a14bb0fc70b21f55de9bc;
mem[461] = 144'hf2391d1002a0fcd1e0b407bb1966f41a0b1c;
mem[462] = 144'he208f8f1ff79fc1bf8ba11e9fd75e5a1e3b3;
mem[463] = 144'hfe19073efd361717ffe6f700edf9f9fa0d86;
mem[464] = 144'hf470ff54f548ebf8f3fa144d056de6e9fcc9;
mem[465] = 144'hee5708f71188fdd4f05ff0e7fc6af8750779;
mem[466] = 144'h1c0cec7e1889e098186d00c31cfaf5fae1b2;
mem[467] = 144'h0b04e5bf1bd412840b85180b05c71a6f11c3;
mem[468] = 144'h1846fafbef25fb63e7dc167ef13cf84aed32;
mem[469] = 144'h1cbd17f9069c17491463ec79f2df1e17f42c;
mem[470] = 144'hf7840a90f3d0fd710f6afdcc18dafeccee76;
mem[471] = 144'hf1d8e89300a002d71a4df535fe2ee76f0743;
mem[472] = 144'hf41c0c71f4a4e989e85f021a0a7deb6ef706;
mem[473] = 144'hfd74fc640af209ea0b0de7e90af5f979ffc7;
mem[474] = 144'hffa2eb72040cf598f4aa0addf51eeaf3fc7a;
mem[475] = 144'h0a9b1363eb520bf20ce2f743f4260edcf3b0;
mem[476] = 144'he66cf19118581e3502d5f42f1672fc780b85;
mem[477] = 144'hf6d1f7500331f4750b5de64ae17b05cb1c18;
mem[478] = 144'h06e51e34e3c61c35e7b7f025ee1a13ea098f;
mem[479] = 144'hec6cfee71fab0e72f4781911fb1703bc19bf;
mem[480] = 144'h0d3e046ee6d6f30a1d28e6bbe21e1d841935;
mem[481] = 144'heeaa19c8e2ebeb49e99afa5efdb4f1b7eaca;
mem[482] = 144'h1e5ef529f554ec4f1c4af814f70be5070887;
mem[483] = 144'he748006e075807761bd41e51e7151063f6de;
mem[484] = 144'h175deda01bbf02f91a940b031124e89c02df;
mem[485] = 144'h0992ee6304ecf07c1d44108fe42ced7ce901;
mem[486] = 144'h0004e3b8e489e752122cfd9710e7ff27f6c8;
mem[487] = 144'h0166e5d9fa5de80713d911afe8731fb1e9e2;
mem[488] = 144'h01051c7cfe9706851ea8ebb10de4ee0f10d5;
mem[489] = 144'he36e0cb304661a02e4ce1a94fd9f1efafbe6;
mem[490] = 144'he5b3197b0d6de934ff14e8f81ced1bd3e057;
mem[491] = 144'h015915471a73070fe5ae13f6e081f285f114;
mem[492] = 144'hf1a01de7f6b60d48f72ee7a3eab70451f617;
mem[493] = 144'hed48e675f494f67c19e4034cfbedf444e790;
mem[494] = 144'h0c66e8bb1dab02e407081a920df70c0e0ffc;
mem[495] = 144'h0ad50f7d119e19cd16200c1ef2ec109201a7;
mem[496] = 144'hfc6b1d39eff113df1dfee924158ff4d81021;
mem[497] = 144'h1255f7b20ad41676f3fe032af7a8f0d40583;
mem[498] = 144'h06db092412f200791cbc18901591f358042d;
mem[499] = 144'h1d74e4e50aca0bef08bb0e540901eac9e19f;
mem[500] = 144'hf6e010a50d05e592ebab131b1d15f4061d48;
mem[501] = 144'hecb6eeff0b0c0080e30deb010cd019f90ffe;
mem[502] = 144'hea16178f0997f26902471a331887f2a90f10;
mem[503] = 144'hf523fed5f26be112f49f14fb161209d9fd10;
mem[504] = 144'hf617fcdee6bb14850afe1efaed2a12ba0d70;
mem[505] = 144'he2ff1d51e53f136207b4f49de9e5efc5ec13;
mem[506] = 144'h1b820be2f3f2f0f9e554fd7d1a3904d5f005;
mem[507] = 144'h130b1374f7d30003e2f9e5110ebefdd0f31a;
mem[508] = 144'h0e0f16b4fb77f3d1085ef3b1f8390458095a;
mem[509] = 144'h16641320e398ec50eff7f3eb1de3f2ca184e;
mem[510] = 144'hf316ff16ff7e0be3fb5de5b5f7fbe22f1e7c;
mem[511] = 144'hf0f70d00f2c019ba1095ec4be7c3e284e4ac;
mem[512] = 144'h1fc91c2ce838f9c7e373e5730a290385ea9d;
mem[513] = 144'h03370edff8351670f3ba115ce7ba0f6310d7;
mem[514] = 144'h1d47ede91381e18de6d0efbbe2a3f336f75b;
mem[515] = 144'he7a4eaa8fafe0ca2098407dde49c1db21558;
mem[516] = 144'he8b9092c0b3e05b005cfe66ee7881984ebf8;
mem[517] = 144'he5471b98f86dff0eea9d171cf429ea06f444;
mem[518] = 144'hfca3043c165afa28edabea34f4d7ebc201af;
mem[519] = 144'hf19b1b770e3c04c30a11e3951d3c089602e8;
mem[520] = 144'h0394f1571e5df87c181c0c4c14bc00300601;
mem[521] = 144'hf099079c1d2d0df60687e12ae4f6e021177a;
mem[522] = 144'h178b0e2709180ac7f9a3e1741d3cf3a3ff28;
mem[523] = 144'hf9ba0b4119b2051917cdf23ce8571dadedc3;
mem[524] = 144'hf7231a950fec129ff74ef913e4ec1a1d0d09;
mem[525] = 144'h1782ee4c08a5ebaef80aefda0ff0f6120d04;
mem[526] = 144'hf9e20447fff1ec60107403c0f7ddfab9e623;
mem[527] = 144'hf0a7ebddeb1a0a440b91f1df08e70c9afd5e;
mem[528] = 144'hedece0d10f5300cd195a0d3b1b0a179415c5;
mem[529] = 144'h16ecff1fe0131f60199cfda4ea0a197ff4c4;
mem[530] = 144'hf529e4ece3360334e3b5ea7ffb20e17cfaf9;
mem[531] = 144'hff840fda0cfa1ba6f87c15e4f76af649f73e;
mem[532] = 144'h139215bdf931fa1b13fe0173e19811f8114b;
mem[533] = 144'hf776099de277e2ad1566153d121bfe57e260;
mem[534] = 144'h1a8bf3e6e680e492f88b12d10e48ef050d69;
mem[535] = 144'hf7ddfc9a0ed6f9e3e707f391ec8e177316c3;
mem[536] = 144'h0da4127b1119ff4be375f2970be0f44af465;
mem[537] = 144'he9c7e29b14900c6a0b9c1b3cfd460ae0e5e9;
mem[538] = 144'h0c1ef909fafd02c9eb0ff759ef66e7e50818;
mem[539] = 144'h1d7502e3f0d60c1d1d080d87e7e8e01d0263;
mem[540] = 144'hf8ad1f47fa12f3f1e52ceae91be00b9fff4f;
mem[541] = 144'h0396e3210c40ed71f581180501320b931b9e;
mem[542] = 144'he0b905e2051c0bc5e1cff1c9e9e212a2f2e1;
mem[543] = 144'hfb40ffabeb0417aff93017670cda0f130858;
mem[544] = 144'hf6fe02e4018b1d13ee9e161c1bfbfb41ea3e;
mem[545] = 144'hf6ae1c6f0e271656f396f6741a471a49e4af;
mem[546] = 144'h19ae1ec2f9c3f1adea7a0a27e4d7eb45fd95;
mem[547] = 144'hf720f56afe20e7b1e1c9f832f263064e1278;
mem[548] = 144'h0b98ed4d09710734f0b7e3c2fb03ec5b1598;
mem[549] = 144'h1f00f1f2e5aaf9e2e0a40fefeb911be30e61;
mem[550] = 144'he5aee69ef5e9f902067c0b0efda5ff36ffb9;
mem[551] = 144'h1f20f3e3fe0b1abf14f214930f37f1abef44;
mem[552] = 144'hf717fad918c9f0afff730ae90e9fe4b903ef;
mem[553] = 144'h095611e0e3a106651e7809a3f998f12110b5;
mem[554] = 144'hf47d14c00875f43ef4b9f551ed6c0cacf1cc;
mem[555] = 144'hfcc0feb3ee5be1ba1d9506b81b53017808e9;
mem[556] = 144'he5f009be0262128ce331105c1e7fef7604c5;
mem[557] = 144'h15d212b7eacdf8e7e3cdedaafba9088cfa76;
mem[558] = 144'h00e8f92ef4741f3a1f9009e9ea61f4501459;
mem[559] = 144'hf547e45206651bdf0513f473ec1af326f8f5;
mem[560] = 144'h1c67ec3ce60ee00a09b9f395e16605aae59c;
mem[561] = 144'hfcc4193efc1ce2be0d0b14a1ee64fdcb01eb;
mem[562] = 144'he006ed3c1dc60c8f01c2f05cf4161719f420;
mem[563] = 144'hfe15f386fa2b06d705f519840f740ecf184c;
mem[564] = 144'hfb9cfc0efcc1e2951f171413e41feb221a22;
mem[565] = 144'hf1efe78a1f74f83d0a1a0e2ae18fe8b10bb6;
mem[566] = 144'hf7d1e368ed8c10f513c11ad10f5c0a8812d2;
mem[567] = 144'h1037efa1f71ae7720499014ce38f0aa0f724;
mem[568] = 144'head5071d0b03ed8aff3b04bd0fc20f67edd2;
mem[569] = 144'hec3a063b1d5f093e02dafbbe193b0437e04e;
mem[570] = 144'hf2d207e1ef791642f8c71b56002f1d6bf511;
mem[571] = 144'h0c99f404fb0deddfe8161f3200f219ab1e02;
mem[572] = 144'h1d8af209eb9119280a07e8dd0f281d94eaf3;
mem[573] = 144'h02da0d5702381d42e967e46e1affe870e7a4;
mem[574] = 144'h09481688f440e4e5f309f85ff8d5e5391b3c;
mem[575] = 144'hee3df15c158b00bd17b2107b09351b070e7e;
mem[576] = 144'h0752ff1c04afe0b20d50f3fbe5b00b6b0b1e;
mem[577] = 144'h0f92eaa018d20280e9c1146d09fe1010e016;
mem[578] = 144'hfeee1eeefa851868e477ea161c8b09fbee71;
mem[579] = 144'he3c314691f46ff5a0ece127be44a17bc0b4c;
mem[580] = 144'h1c9e0edb1f5ce312fc3ef620e80a192c085d;
mem[581] = 144'hee900d59f0d7eab5168f017b11b1122600ad;
mem[582] = 144'he35c1e16e5d71bd4e61603f403ece2b1ed3a;
mem[583] = 144'hfc8b1c2e15c8035ff17c0f1a00eee4c9fcdb;
mem[584] = 144'h099deb851499055a053d1454020a1d6bea18;
mem[585] = 144'h11defe020c32f831f4e30fcf029b1095e4f1;
mem[586] = 144'h0676153910dcf8f61158f45e0235e351e73d;
mem[587] = 144'he383ff0e062be8bd0f2d0eb0e9c21a28e9fa;
mem[588] = 144'h08abfcdef58fe0111bec1d3103140579f678;
mem[589] = 144'hfef805871ea2eeeaf1f10a63f44e0dfde9c3;
mem[590] = 144'h14fbe043ee7b00ebe947fc1fee66ee030f70;
mem[591] = 144'h1fbc1fbf12f1eb7af3c5ecd3fc3605c20637;
mem[592] = 144'h0a7be157096cec6cfa1feee2ebf2e2370a3e;
mem[593] = 144'hfd34165c044d0a5ae514f3d3189e07460926;
mem[594] = 144'he9700712f52de196e0a7f1b416b116d4e774;
mem[595] = 144'hf51f1edbff1001e809d11a2c1076f55a02ea;
mem[596] = 144'h1ce0e6b4e5fefd46ee6b150de5ea115405fe;
mem[597] = 144'he8b304f1e2fd1743f8361a50fa6f0a481352;
mem[598] = 144'h14a2e602f0911c3e1114ece4fa561cbe1cd0;
mem[599] = 144'h1622f5f8eac3efe6e61afa87e79ee377197d;
mem[600] = 144'hf59eefd5ee3413f61a5ef008e2a3e1da0241;
mem[601] = 144'hee6def28ef0f0764092ce3f1f074eadee861;
mem[602] = 144'hf0d4e56efebdee17fc0808a0e2f00d6b1157;
mem[603] = 144'h008cfbd0ec3d0b301e840def18dfe2d11ba6;
mem[604] = 144'h131be4d5faeae78c1b62068511611953fd00;
mem[605] = 144'h08c5fad1f464fffae8a6113cf51e04560118;
mem[606] = 144'hfae208aae96ee43b1dbce301158be95f047b;
mem[607] = 144'h149e1de016f90c80067019cee6c9e73a102c;
mem[608] = 144'hfe460ad41c510265ed63fdb219d2e6060472;
mem[609] = 144'hfd87157a192e0e1b09611890f55607a8f67f;
mem[610] = 144'hf429efde08baf5d6e5def31eeb1bf156e892;
mem[611] = 144'hf0ee1e03e781ee33e3f7faf8ef68fda21987;
mem[612] = 144'he20efc74fdfa1473ebd20e66eee412b21172;
mem[613] = 144'h19b5e8210ed708ec0da2f1c0fec20ed41949;
mem[614] = 144'h138609f2ececf3cb17e6f054e3defc8009b8;
mem[615] = 144'h00171795f78beb2fee64eef00920176ff188;
mem[616] = 144'h017718c413a2fbad103aeef5fdb5eceaf365;
mem[617] = 144'hfd59fe9600c6e4b80cdbede1fffb1c651baa;
mem[618] = 144'hf3b5e1a8f5e9e58e0c380eb7e2a5178bfdf4;
mem[619] = 144'h089b0433e486fab5f7760ac5f975fe341c17;
mem[620] = 144'h0a04031c049eeda1f9fb19db0df0ee750546;
mem[621] = 144'h12b10f25e631e9eb19faf5edfa501f350b5d;
mem[622] = 144'h031d0c8202390b590018021916050f32e286;
mem[623] = 144'hf826e146170611701895f5b50edef8c0e3f2;
mem[624] = 144'hfc30e2f2e4ea163e169cf866170910c10e84;
mem[625] = 144'he5aefe25015907330f1be342fd6a06e3f093;
mem[626] = 144'heaf8012716f2fafb06e1e061024c19591ca0;
mem[627] = 144'hefbd04e816eb0fe2e9cce486eec8eaafe663;
mem[628] = 144'hf1adff650c650cba0cb0f596ed84edabf17a;
mem[629] = 144'hfb94ea9cf6e5016af8c4e6d7efcfeb531f03;
mem[630] = 144'h15f5f7bb074a0956152207d20009fb35efa1;
mem[631] = 144'h03521b9107a31b71e8d8e949ea6d18c7f4be;
mem[632] = 144'h07dde8b9f0a1003c18b9f1400c4fea6f06e3;
mem[633] = 144'hf0ab102d1cdbed65f8921052eeb0fbe6116e;
mem[634] = 144'hf28be0b0e8aae7fc1f90ed7410db0f86067d;
mem[635] = 144'hf309f0890a36e79200a9062df24ee8821fd9;
mem[636] = 144'h16c0ed6dea2ef63b121be404f374fb601d19;
mem[637] = 144'h136f11d4ef77fae6e7f7f413e07413baf73f;
mem[638] = 144'hf18019620ea0f65c1e980e9014e90c631357;
mem[639] = 144'hfd99037a14f9e6ed1d140788eaf3fec7fe70;
mem[640] = 144'hfb7deb920399e0521279ecbd039909a21026;
mem[641] = 144'he07017d7092a1805f2d60f6a1682f630e5bb;
mem[642] = 144'h05f20d9e1271e51ee396eea2f2dfed58ff81;
mem[643] = 144'h1ca7eef1f5e2f085105a1a14e0c4fdd7e5d1;
mem[644] = 144'he4560c711c4703321803ed890707ec60e087;
mem[645] = 144'h03e90e3210cf0dae1b5bf6adf7dbf7c3fa02;
mem[646] = 144'h0a5e03c218ee1acc1ab0f81101000fc6f17a;
mem[647] = 144'h0f89f595ec42e7dcec04f1d2e3f01ebd0dba;
mem[648] = 144'h0b7cf2320fc80b21eb2aedb71315ed17fe92;
mem[649] = 144'h1106f6201e1ef408199dee8deaaee3590304;
mem[650] = 144'h197a13950876f142e6bdf894fdf61df40331;
mem[651] = 144'hffcce6f8114d0c41f426ee41f7fc0863ff32;
mem[652] = 144'h18db01d1f298e39001e1e3fdf19a1b7a0ddb;
mem[653] = 144'hfb8feb71fae71697103ffb9aee2414501713;
mem[654] = 144'h09e408dd03b508a8163002fc10bd1169fcf9;
mem[655] = 144'he13f1bda088ee163192e1ccdeccc1d0e130c;
mem[656] = 144'he6cdf6a41bcb1742ee890decef8cea5ae4a5;
mem[657] = 144'h0b6515aae66b11471356fcee189f030a0815;
mem[658] = 144'h0a16f0a20276e5140a1e0ae319c91db50fe3;
mem[659] = 144'he214f2b2f440ecbeffbc0737e87bfd35e231;
mem[660] = 144'h14ed1b92086becdc1137f5c0f9400964f12e;
mem[661] = 144'he0ece1c61214e51efddbe76915c90d21eedc;
mem[662] = 144'h1d8216530ddc0941fa30f6f9011eef93e622;
mem[663] = 144'hf16ff15cfd5d133ce9c9f20203bd196e04a3;
mem[664] = 144'h1b15eef9f93d1098e4bc1e30fd83f3f40435;
mem[665] = 144'h156f19ee11691841e58d1654f452f9c6130e;
mem[666] = 144'h1abee636fd4e1527ff2be7820b831c310c0a;
mem[667] = 144'h17391dae093408b0e816eba5f3ab18d4002c;
mem[668] = 144'hf34916db1a3912731d34f7e0eb40072b0fd8;
mem[669] = 144'h0c08019bf005e050e4411d21ebf0fafcf677;
mem[670] = 144'he4fc0c65e6fcf76f1fcce7c0137f171a1bb5;
mem[671] = 144'hf43409ac1302fa77f2a3fb1f0f35ea9df9b6;
mem[672] = 144'h02871823e124eae2f16b12d318601cfe08fd;
mem[673] = 144'hebbdf2b6fb5a1eb70a3b1154035ce875091a;
mem[674] = 144'hf655e7570f78e4a204da1ed4e535fa85f3e6;
mem[675] = 144'h19fe0b1ff82917c7f89a1006ed67e82ef4bf;
mem[676] = 144'hf95de9ee077f08d5f0bbfd650e82e71f022b;
mem[677] = 144'hfe8ff107e1d01b5f019106c81859fa75e8ca;
mem[678] = 144'h064312f21760ebbe188be1d500670f8b0b8b;
mem[679] = 144'hf8ba01ac0fa8f5c0f1c9fac6e93ee82e138e;
mem[680] = 144'he58df10ae0b7011cf13c1c6ae53a170ce90b;
mem[681] = 144'hf35509d3e331ecffe26ceb76069f173c0421;
mem[682] = 144'h0118f56fe2310a5713f0e842062eeb06013d;
mem[683] = 144'hfa35e46e085e11d01456e2fd125111251890;
mem[684] = 144'h0de3fd951129e5330eacf83c0afc170b0a81;
mem[685] = 144'hf34ceadcef15e643e4e91b41ec901b2ee971;
mem[686] = 144'h0c2a164018dee66f0a111cb21846f23113ae;
mem[687] = 144'he2fb110b0c39076a01b7e5800dcafe1ffed9;
mem[688] = 144'h17cfef84110ee4671a7201e3094ef61ce8c8;
mem[689] = 144'hfc4de341e1e3ed34fea70d5c13f51115f4ed;
mem[690] = 144'he370032d0f56199de4baf0651265eeafe07b;
mem[691] = 144'hf79504b817ace1bdf2730523edb508f3ea9c;
mem[692] = 144'h0532e35f0930e2e71f1601d71d860061ee69;
mem[693] = 144'h15611d85133ae1a6e1a8f6d3ef7eefc8fbe9;
mem[694] = 144'h18370e46158e164cfe8f111dfb07f22b1b75;
mem[695] = 144'h103b064d1338e6a50af1e208f791e9e30430;
mem[696] = 144'h00bee129ea5608f9ed9419190b930085fde8;
mem[697] = 144'hf9f601ad0157f063f09ef299fe32e33519a1;
mem[698] = 144'hffaafa4e00c51c2fe46f0bc201d80d7ae937;
mem[699] = 144'hfedc1fd8fe6119e60fa207a90f44e72f0c5a;
mem[700] = 144'hf4b3ec29e3fbeadf1af20a65ea56f6dee033;
mem[701] = 144'he013e095130c1baff266e7cdf1e6f0ee1ac2;
mem[702] = 144'hf4fe0321ec30edd3fcc7101ee83c054b1c8f;
mem[703] = 144'h143ce56f1bf10ceaf0f8f030eb11ef221fe2;
mem[704] = 144'h143e196d1ca0152ae3c3e17bf3741e1b0e21;
mem[705] = 144'h138be3f50d7d1f4f05d40f2e0d4109d6e364;
mem[706] = 144'he305ee02fc761e09ef7507a0eb29145c0766;
mem[707] = 144'h0a67ecc80203e253ebed1fa619f8195f1fe0;
mem[708] = 144'hf5fc06f5e9b30e21e2d4f9ad10040bd61a66;
mem[709] = 144'he3b4e18c1a3aee0bee0a04ce0c99186e158f;
mem[710] = 144'he35b0486e1231e9ce201ef3109ebe3db048f;
mem[711] = 144'hff95041b0bebf6c1e6d4fb52ece013f816b3;
mem[712] = 144'h0631e6bdead1e722f509e22b149505b6f9d6;
mem[713] = 144'h1ba9054804ea153cf4be1f8111a8e32215e0;
mem[714] = 144'h185a1f78e0231caa083a0d851d3605a5f7f2;
mem[715] = 144'h13221c0111cf09f90622ff6efd69e36ce7c4;
mem[716] = 144'hf23be5bc1f771099121c061ff265033c0267;
mem[717] = 144'he08b1bff14fbf292ee5bf58a0e681c721e01;
mem[718] = 144'hfecd048a13451e3aeeb8f322195bf22e126d;
mem[719] = 144'hf46e133ee0c71dd515c81038ec8ceb11f034;
mem[720] = 144'hfd9e184213c0f30d1318efe5fe01e3b2f233;
mem[721] = 144'h0f4eec410b17f34205f115cffb2002f40f1c;
mem[722] = 144'he393f3fc1672f90df67a1e330e15f714f6e9;
mem[723] = 144'h1d081d54e19dfc091ca5ea9ff1c7fb5efa9c;
mem[724] = 144'h1e28ef8cefa9fb28f606101fe50aea0de737;
mem[725] = 144'hf48312fc1d5e00aa14090781f12f0c5b0b90;
mem[726] = 144'he17cf8a7f566f4cf1d440a9e0e2307361a9c;
mem[727] = 144'h0a93e7faf6ad176cff9ee36ce0080155fe71;
mem[728] = 144'h0f540946fdfaed920a51f3351c69050afccf;
mem[729] = 144'hece306080f3efc380f20f99a148ef3cb1582;
mem[730] = 144'h07721ed4e11ffbed18baf9e6f9def7abed2a;
mem[731] = 144'he34402e3e3c5f94204ef06eb1353f2c50ee6;
mem[732] = 144'hef73fa7a08afec260477056efc50031aea30;
mem[733] = 144'h1bd2e9c906531eb4f923fbf8f3e71d59ea50;
mem[734] = 144'h0a3a06cf044a08d1ee65f151f926ff441744;
mem[735] = 144'h03bbf86fe9b10d0c0657134e163806ac173f;
mem[736] = 144'h00f80d2a1749efbe157d136af568ea9d148b;
mem[737] = 144'h0a20196615d61fc40940157be49013801ffa;
mem[738] = 144'he4941e48ffa6f412e81cff80eed900190986;
mem[739] = 144'he606f584efe5e434f97a0d5de637eb411047;
mem[740] = 144'h069e03bb033601030b15e1b9178df7e5f10c;
mem[741] = 144'hf8b1122e1bcfe8f8e6fa0e20fc360b7bf361;
mem[742] = 144'hed221821e397f04703630fe70aa0f83a08d3;
mem[743] = 144'h19b8044a0235f70ee4051c0113d712b21205;
mem[744] = 144'heb270c93f842fef9febbf5f1e72cfdc60c63;
mem[745] = 144'h11300901150f1cc119581c16f1fefc46ecab;
mem[746] = 144'he946ee0105fd00f6156ce06a13a00049e1f3;
mem[747] = 144'h00f51694e232f85bf0b21933011316151472;
mem[748] = 144'h1555ee591f1fe924e81cf7f405ed0fbcff50;
mem[749] = 144'he7601e69e9a9fdfa02690cf5ed51f2e91f34;
mem[750] = 144'h00740b0cefa1f1aa1befea80ee71e2f21e6a;
mem[751] = 144'h012fe36301fef9d21662ff6018e307d30a13;
mem[752] = 144'hfd37e9d3e0d1fa62f6391181f737e1970f23;
mem[753] = 144'h1c9a052517f2047b00d4e29fe770e7620518;
mem[754] = 144'he101f3ca1caf03690f52f344ed420fda1624;
mem[755] = 144'h0bdce9940e511eaee8e8eaab121af2e00c5f;
mem[756] = 144'h0abb0b6def721a52e3a2f7faf73813bcfeb5;
mem[757] = 144'h0e84e63818b5f025fc3403aae629e1fcf7d1;
mem[758] = 144'h04f90fc70b0d0464f22e0e9fff9814661e37;
mem[759] = 144'hf565fe43f3421ba702301c6419cc06f01fa4;
mem[760] = 144'h03601f78ed5e083bed8bedb51babe47befbc;
mem[761] = 144'h0846e84509b905c60f811f410a14faca0965;
mem[762] = 144'he71df7af0d81e3aaf687f6391fe01544ee6e;
mem[763] = 144'h079a0687e249edf9e41f17c9e3f70c030b58;
mem[764] = 144'h01fa1a571c711081024c02b7e66a06dfe19f;
mem[765] = 144'hf04affee009d1ae9ff72e427ec701da3e6aa;
mem[766] = 144'hf0eff5a6f56bf0bf05411777ff8b07e2fad5;
mem[767] = 144'h1dbf12c11ca11d50f8a0f4bbf0580da01b6f;
mem[768] = 144'hec721f55f9870537e93b194810820bde0932;
mem[769] = 144'he940180b084df8e01462159ff9d5e85905c3;
mem[770] = 144'h1e511c8f130f12b1fc860637edd5153de67d;
mem[771] = 144'hfa65f504fbac084002a6e5140ab9e3c21152;
mem[772] = 144'h1741fddb00430ffae37eebf313021a320a4d;
mem[773] = 144'h1de70db815831a1f0b4cfcc5f3240964eb65;
mem[774] = 144'h115ce454ef3d0ee9f98b141de627e33f08ca;
mem[775] = 144'hf2ebf1431e8f102f032a0494fc3411190314;
mem[776] = 144'h0c541767e8cc178b15311efc0eb8ecb4eee8;
mem[777] = 144'hefdef206f96b02df01a3f291e7d0fd1fe4b4;
mem[778] = 144'he970ec48eeeb17b1ea7b04bc080dee18efb6;
mem[779] = 144'h0814fb9ae828f787fbf51b32183c1bfaf009;
mem[780] = 144'hfb06e38de8d7eb76001cfd9f0f54004de99a;
mem[781] = 144'h17bd1c48eb761869f0ffe28c07dd19b009d3;
mem[782] = 144'h01deeda20ca900670b20e52301231a2be11a;
mem[783] = 144'hfe43e962f043f1bf0918ffef189f1d4bf869;
mem[784] = 144'h1715e4b50a831aabe4eef3fbe242012a1ac1;
mem[785] = 144'h0c80fc70f6b0ff89e129e441e158123615a6;
mem[786] = 144'h0f07fa47e8841318e12102c71e82f93f05a7;
mem[787] = 144'he728e73df0bc0a01e1f408950736e3da1a63;
mem[788] = 144'hfae30a2313481d930427f7cf1254ea491580;
mem[789] = 144'h1e18e2fa1a4a026cfd7af61d1db3e39af6f6;
mem[790] = 144'h17d0e2a4fe650847f4790f5e13d7187f1341;
mem[791] = 144'h078f1ef9fc550936157c1150f76a1c3efd2b;
mem[792] = 144'he180e2750c17eb01ee24f39af37ff99ce81b;
mem[793] = 144'hf8d11672f81b0afa1d8219a21077ec3b1957;
mem[794] = 144'h1db4eb73113cf499028f0214f0051d3eeb78;
mem[795] = 144'h0227e3b80333f745035cf9b1f0bcf2c11704;
mem[796] = 144'hfa77003c0e191c07ec891613e84be6f41aec;
mem[797] = 144'hfa7c11f6007bfae91c1fe526f70ded110212;
mem[798] = 144'h0875f61214bc04630d0e1a7beff00eabecfb;
mem[799] = 144'he5470d1d07750edefbe0f9edf07c07170416;
mem[800] = 144'he11eeee1e8441407132fe3a4198e13c00f2c;
mem[801] = 144'h118213180706ebe41e481ce2f25e1700fc70;
mem[802] = 144'h1027e0a9ef3717400ba1e84ef870e62f0546;
mem[803] = 144'hff7a1167ec1ff4fc031a034bf601e1b5f3e2;
mem[804] = 144'he4b313bc0a77107909a9f52df5350f3b089f;
mem[805] = 144'h0818e3fb043c16a5e148e3dbfaab0f33f015;
mem[806] = 144'he52d1681e37ee1c3122d0940f94fe5251846;
mem[807] = 144'hebaeeda1f2221a1bfd3ff29ef7590a7a1709;
mem[808] = 144'h0d1e0cd60a650cde0e4a0d06026d03dc0333;
mem[809] = 144'hf065ec0ee39ff5c1efdb1553e169e2a30c9a;
mem[810] = 144'hff68078eef85ff97106dee9b17de08fa14d2;
mem[811] = 144'h195af3ee0e75f8650987e647efa2e058f39f;
mem[812] = 144'h14e00fd91e46ed52edeff49411e60010fce1;
mem[813] = 144'h10e50aef0f3d10cdfb44eb850e0410ace06c;
mem[814] = 144'h0df3e536f1a50e500a3704320acc10081a11;
mem[815] = 144'hf2351c96fe0f1a17e90a0337fbfdee5719ff;
mem[816] = 144'hf5e41f4f1d0402851f8bf849ecbb1f0d0bc7;
mem[817] = 144'he66df44d1c32ebfe0062f90f0b3fe9620b44;
mem[818] = 144'he222f3d8e82d13121860035808a9f0fc0165;
mem[819] = 144'hfd8a12b9edbafe6ff962116d0c2f033bed1a;
mem[820] = 144'h17c516d0e25afc0aef2be12f1ccd039113a3;
mem[821] = 144'h168012821863017d0c31fc6b1b051f02f895;
mem[822] = 144'h1667059115caf2eee05de656f7d115861d3c;
mem[823] = 144'hed94efff0b4bf56509e8e5f9f26d0f1f0f22;
mem[824] = 144'hf82ae665ee7a033f0a56fcf30c13fb93030f;
mem[825] = 144'h1963f445f9a81ef604290a9bfd8f0839ece1;
mem[826] = 144'h08551c5f0ac10688f1d61ebce39e04df0687;
mem[827] = 144'hf852e048e7270ffefbac0d76e0170d9b170b;
mem[828] = 144'h0e2ef7d5e679f23f07940309152e0687fece;
mem[829] = 144'hf194f41bf49efb12f89d128cf9f0fb4c185b;
mem[830] = 144'hebf8e802fde2efec1ef31475e37d1a7bed47;
mem[831] = 144'headd0615115b1489041becf019aaf158ea0b;
mem[832] = 144'hf0e906b6128ce594eeb30a811e811198fb91;
mem[833] = 144'he95be19901d7175ee5d90cc6038409e1ee3d;
mem[834] = 144'he787e9ef022fe069e8f3e98ae2fb12affd18;
mem[835] = 144'h18220593fface10a10b3e383eef30409e4aa;
mem[836] = 144'h0c750d7fed50fd27081f0bdb1506ec0604a3;
mem[837] = 144'hf27b11a2ed7b165fee8cee2308190cf8ec91;
mem[838] = 144'h1b8c0a4e0664e7be0f071ff6f4260c97f3e1;
mem[839] = 144'h139b1cdffe29f9901e6717c61572f013f760;
mem[840] = 144'h1d5313c4f6521bbfee771c39f866fdc6e63b;
mem[841] = 144'hf97611aeed3ffa05064809f3efe712f70856;
mem[842] = 144'hf945ea31e93f0624142aef5aecbefc6b0d45;
mem[843] = 144'hf786102d1976f8b3faad1bbb0c9ff3141fa2;
mem[844] = 144'h064a046efa0a1ea310c41ca01e60168ee7df;
mem[845] = 144'hea17f6851530eca60f23e51f1b91f269e82b;
mem[846] = 144'he5ad1766e4421d8af1761350fbebf42b0733;
mem[847] = 144'h05f1026411f000590e5f06b7021efc70f21f;
mem[848] = 144'he96cf2bdfa6614090d76ef5ce4ec0ebd10eb;
mem[849] = 144'hf717e683f0d70982f4e2f7c2f6f70131f384;
mem[850] = 144'hf0b91f9fe3a11ae013e5f08ceeda1bf61dde;
mem[851] = 144'h0a41e511e21deccdea6be2fcf3b7f37e0595;
mem[852] = 144'h15daf0daf9cd00be01ec0b0808440c29ff78;
mem[853] = 144'hf8271f311249ef3fede90e620cf30fabfca6;
mem[854] = 144'h026805a1f1e3e93206c8fac2fa3c069d06af;
mem[855] = 144'he6f50f8e10240c960e35f6631e75e62d1c19;
mem[856] = 144'h06b2e4820f7505c30f7af8440fc51ad3f485;
mem[857] = 144'h17bd01f9137d1d390ba6efbb0e3803d4e136;
mem[858] = 144'h12a4162f01bff3690fd3fddc1b6e066001f6;
mem[859] = 144'he74e1d0c1e8fe973e350eb5bfa88fac2fb01;
mem[860] = 144'hf428f408ee17fe6ae7391b90f183e054efae;
mem[861] = 144'hf231f57209cd18caf6f2f7891ecde04bf54c;
mem[862] = 144'h138514bef55deb7be61f12391595125016f7;
mem[863] = 144'he8ac151c0185f2aaeeb2e28510d7e30602a7;
mem[864] = 144'h1cd5e614f82b145e0d4c1c15edf4e2f0f857;
mem[865] = 144'hfe32f406fdb61ff40eacf7f4e0d0e059e00c;
mem[866] = 144'h192dfcd1fdfde126f02f01d617fd045febab;
mem[867] = 144'hf1caec59f7d916f2fdf50548f6de104a02b8;
mem[868] = 144'h0b48f2f31ac4eef300ea1550f2ebf330134c;
mem[869] = 144'heebe1c7efb1be833e5ed0fd5037e0528e5f8;
mem[870] = 144'he35ff08d1e2f0f430a9fe4dd00fc0142f1d2;
mem[871] = 144'h0b5900bff2beefd609630a60edb711cd0bba;
mem[872] = 144'hfae6095fe6a01c3d191a18f61c5efd9ceb2e;
mem[873] = 144'he6c6f6f5eb6312d5067fe725167c0d2d13f1;
mem[874] = 144'h0c200f67ed720decfd58088dfce9f3b6f898;
mem[875] = 144'h1cb41e090f22e587ea4705981472f46e1e51;
mem[876] = 144'hea55f2c30757f1980c5609701fa212cb1cda;
mem[877] = 144'hf004fa150b61f6dcf7b9f268e8620197f457;
mem[878] = 144'hf25ee43c11290bce06d61e9cf749f7c5ee0b;
mem[879] = 144'hf6dd1899e801f725e2d60420e865e9e000a5;
mem[880] = 144'hf466e0bbf42e0116f574fbdbe8ff1ddaec42;
mem[881] = 144'h1686e9a8141df00c12d202060d3e0c92f0a4;
mem[882] = 144'h1e3602e51ee4e1e2e190140efd731c0903cd;
mem[883] = 144'h0a0f11a0f6d4e45305fe10c0edde0af30939;
mem[884] = 144'h0ce4ebe506e9fc240ce7fbee077d0877fc3a;
mem[885] = 144'h1ef80ee3081909100267f0b3f86e1ca8f08f;
mem[886] = 144'h18c10b80e58ffd8215880f71f218efdae4ad;
mem[887] = 144'hec79fd1f1090f43ce2c9f6fe0a9f0d3ce3dd;
mem[888] = 144'hf73c09ab142d182b0e2eefa217d9edf4168a;
mem[889] = 144'h0a4f19eaf8681cb3f3631d01e40dee9ae0e2;
mem[890] = 144'h0d74f89a007a11ce00041fa8121617adff6a;
mem[891] = 144'h1b001498e6e70de812211cffe98b025f183b;
mem[892] = 144'he55be45ae2cae29ee3d4e35b1e4a0c1e1138;
mem[893] = 144'he690eaa51eb31a1c03a1f230fc3517c4e850;
mem[894] = 144'h05890487f89c0ff9ef1212ed0f880249e360;
mem[895] = 144'h010ef73df29815c3f0091c6f1bcfe48009c6;
mem[896] = 144'h15e105edf0afef561605048bf8ed05e0fb36;
mem[897] = 144'h0f63f9ef01101f930adc1f61147310e603a0;
mem[898] = 144'h1f9ff0ca0ba90d8801f70dfce03206390818;
mem[899] = 144'h094ef69ef195f3e3e576ebdb0b581c260645;
mem[900] = 144'h194f065cedf9e93bf7eb08b01f44ef17e321;
mem[901] = 144'he0771d491f8fe6af05dfe03bfd0ae611fe3c;
mem[902] = 144'hea3b194ae2fe0225e5661ffbfe640d12e94b;
mem[903] = 144'hf7cbf3bb0cdf0d3b0636ea8ffc350ce91ac0;
mem[904] = 144'he2630cfdf8e1f7befa4ce6291fc2f14af6a7;
mem[905] = 144'hff02e415f0e5fffef4b113220abce4b91613;
mem[906] = 144'he76ef0ad00381f57ea6815aef0caf565f532;
mem[907] = 144'hfce7e54f0a8f0167e97208bfe4140087fb39;
mem[908] = 144'hea24f624e4bc10470e66e8bd0ef911b4ffab;
mem[909] = 144'hf392eb6ee252ff371c89f0ef0e60ee2c1b03;
mem[910] = 144'he468fa37095aeae018b500e3e2d5ffdb044c;
mem[911] = 144'h1dd1e58bfbcaef20e2f0fc52002b1ae602e1;
mem[912] = 144'h0a25e3f6067a0708e051fe1c0d921e680e22;
mem[913] = 144'hf2ab13aafcdc1243fac6f1a2e32e004f10c5;
mem[914] = 144'hf632187a17b902741bd4000dfdc11f2fe1e8;
mem[915] = 144'h196c15b1f0ea14e7ffcc024b0f1bff0bfcca;
mem[916] = 144'h059811d0f655017f074c0a91f604ff511f33;
mem[917] = 144'h0c61e84ce8e7f147e38411c51a111a7efb34;
mem[918] = 144'h12edf8520732f2080c600322e1d402d2f474;
mem[919] = 144'h028a0d9c05770180ff590739fa69ee62eb6e;
mem[920] = 144'heb29fe4af333fc270db6edaaeeb1e0740190;
mem[921] = 144'he6dd1168e142e718ea17f0960b47f97fea2f;
mem[922] = 144'h1be4123001d3fedf1dbaffed1f48f3f008bb;
mem[923] = 144'hef82f6ed14e4100219fe182b04470ea21b66;
mem[924] = 144'h11d91f2b1ac1ef38efe41efa0b04f0cdf54a;
mem[925] = 144'hf8f7f768f519e1660a0c1b77fb7af923f438;
mem[926] = 144'h028e0708f2d61a2ce8e1ec24e339f83a114b;
mem[927] = 144'hee80e32ae0a105830b3010d90fc4e92216b0;
mem[928] = 144'hf56b1e90e626f105031417fde216ec3d1e1e;
mem[929] = 144'h0e00fa91ebd9028ae3341651f7851a3ae4bd;
mem[930] = 144'hf2b5e698ffc10192113c193714bd10c90917;
mem[931] = 144'h1878e8910fa6072911b804b7e0a40128ea66;
mem[932] = 144'hf4d0e621f126f9d8f3abf6c5ef5610870ff4;
mem[933] = 144'hf8450a9cf6fee5b6eb8c1f2b0b73ff6ae1b6;
mem[934] = 144'hf3a8f3f91dde15cff5f305f6e8e218ac0346;
mem[935] = 144'hf0121a04f2511eb0eba9e533162c1abffd87;
mem[936] = 144'hf9c0e7701686ee651c42fd9ee9711491f55c;
mem[937] = 144'h0a4cefd1055603e00637000ae260f3e50d24;
mem[938] = 144'hf4a4f4bc1416020fe5ececa8066e10821b39;
mem[939] = 144'h0070f0d8111c028d05d9e181f66df294e39d;
mem[940] = 144'he20ce8a809c01a0be210f5ee0fe7fd3513ed;
mem[941] = 144'h0d3bfedde8bff78108b10cd4e85b07ac10f9;
mem[942] = 144'h197912a5fb45efc219b8edaafb3c165a10bd;
mem[943] = 144'h0c51fd9af50310651736fb65edc9f723e3ba;
mem[944] = 144'he2580d4f116feeace54016a109951b7deef9;
mem[945] = 144'h03630398eca3f85117f2e2bee057e9bdea8c;
mem[946] = 144'hebfc14b5f2690025f9e71cd917cdebe015a4;
mem[947] = 144'hf5730caee86d1a89e89006b7f6c7128210f4;
mem[948] = 144'h1facfa3df8aae385e5f2f463e00607b10509;
mem[949] = 144'h0db0f850e0faf21dfa3106cce781f51ee958;
mem[950] = 144'h09c2ea0ae7fbea10102be9e2e797e84eeb57;
mem[951] = 144'h0e06fc71e591f75a19331ca90020fdc4f713;
mem[952] = 144'hef5b12dc047fff881bd913def8d11b5118fd;
mem[953] = 144'he4641710eee008f804f4e358fd35f024f7cc;
mem[954] = 144'h1e82f83f11ce0b7c1aa0e289fae1f08e08b4;
mem[955] = 144'h1842e9be1ba2088418b2e5500fcc09d80df8;
mem[956] = 144'h170408cc0775fd7c078af8d7095614d6ea46;
mem[957] = 144'hf10607cff5f90a2c0b1bf2810f44e3b2e3cd;
mem[958] = 144'hfa54ec9a06b703b5e18fee66154bf0a0f42e;
mem[959] = 144'hf963e1fffa0007cae2410546eb3819431fc8;
mem[960] = 144'h0060f28a0822f170edc0f1e5ff6e025113ac;
mem[961] = 144'h03ef0bf0fe601980fbf100131936ee38e838;
mem[962] = 144'h0f90fb57ebb6e4340df1fd97f3450112f94a;
mem[963] = 144'hfb54ec2e136618950cd0e29cef5b048e1eee;
mem[964] = 144'hed4808661836f7510a6d0c251a32efdcf563;
mem[965] = 144'he82c027e00f81a5aeab8f700f7ac16eb0a4f;
mem[966] = 144'h17f40af0f7c4e177e86808bf00b4179a0394;
mem[967] = 144'hf48e1190ee5107aae9cc0807eea7041cfeb9;
mem[968] = 144'he8171404f66d14d504440903e4dfffcce76a;
mem[969] = 144'h0dfef5880a5109dd1445fa7ce7c4e86a046e;
mem[970] = 144'h00f01ce906a7e557e70a04e01bd6e85907d9;
mem[971] = 144'hfa8d0b121d211231e36e0f5f19f20360f818;
mem[972] = 144'hea04ff620a740e3601370c291d19fc27ecc7;
mem[973] = 144'h1e451792e293f88efe1be7c316c6ec31e7b2;
mem[974] = 144'hf97cf3701b3be64800eb1fbafbe2e9c3f4ef;
mem[975] = 144'hfcc11940f0dd1e3812ade5780d6e0a41088e;
mem[976] = 144'h06fe005d168a0e4c1a26fc2f1dfc1940089c;
mem[977] = 144'h1d221708e46cf991e5d1158615abe0980216;
mem[978] = 144'h0df41ae71d85eeb9fecef268ef1b08f8fbfd;
mem[979] = 144'h1371f965f37befb3152bf14a1b5e110ee929;
mem[980] = 144'hf25210fb0386e64fe1d4e1af082a09ce05f9;
mem[981] = 144'he4f71bfd078900ef18821db71640e1b00593;
mem[982] = 144'he94e0208f184065c0e2302f31c171ec70a8a;
mem[983] = 144'he269045b17971857fd64f1e50d9208c2e17e;
mem[984] = 144'hfb77088c0151ea78e24303bf00d50a2215aa;
mem[985] = 144'h03271acde265131bede4f1c8fcc703441d22;
mem[986] = 144'h00c8fc251ba0e6ec110beef0f77004fe0edb;
mem[987] = 144'h0dcbe2bced87e803fdd81487e573feb9e843;
mem[988] = 144'hf6cd05161cf2e3c4e0c6fe89e9c0e3f7fd8d;
mem[989] = 144'hfdd3ec96f02cec68001cf02716daeacaebb9;
mem[990] = 144'h10d3ef061f29e88aff9719961b3c00520ba7;
mem[991] = 144'hfe69feace441edfe1df3eab51ad50814fa82;
mem[992] = 144'h0a9512b51967ee481a40f66d1bc110cde34c;
mem[993] = 144'hf73d15e8e7c0e2df1e4b01cde27d13e31223;
mem[994] = 144'hec1701ca105fe77dfc3c1b4a1538179ae55f;
mem[995] = 144'h1b14f5b1f5f11d5300d7eb7310d41ae314f3;
mem[996] = 144'h15520100f4cb070af89c1c281252f52b19b4;
mem[997] = 144'h045e192ae939f0771a0917d4f195edadeb86;
mem[998] = 144'h17a313dfe8270973e198f234f6d3f7b4028c;
mem[999] = 144'h13f5e6bbeccc02081cd9fff8fba70bf4ea68;
mem[1000] = 144'h1f43f4a4f4181a3de3d50b80e4c7f355f171;
mem[1001] = 144'h1efef7b7ea601472eb0af18019c3f43707dd;
mem[1002] = 144'he78cffb109e1fb22ff4afba6057de87d0544;
mem[1003] = 144'hfbe8e26f0c130603e71af1cbfd62f186f28f;
mem[1004] = 144'he03b06cef07ce09e163c01cfea0e10c81d14;
mem[1005] = 144'hf8ed164b057b00a0f40a0aa50638fd0c1c89;
mem[1006] = 144'h13ea16be11490a5317c1164ce94d135ff04e;
mem[1007] = 144'h0bdbfb8be4181f2a16a20351e33d1d460746;
mem[1008] = 144'he59516ab09e4f8d3e359e593f2fee67416c5;
mem[1009] = 144'he6cbf989e1e1e27befdf19e011aa1bcde1b9;
mem[1010] = 144'hfbc617bc1cd31f581c50ffc4fc0406680535;
mem[1011] = 144'h17781b0d0a33fcf2e04f01c6f848ed761864;
mem[1012] = 144'h114ce2ff0982ee4ce49c08190febe7a115f3;
mem[1013] = 144'h194cee62e6def5c8fb6afbd6fc06ff05f633;
mem[1014] = 144'h173000f5f8b2ff4bf9e50a181c4dec701832;
mem[1015] = 144'he2e6f9f2e22ee7fb05f10cc1fa9fe49b11d3;
mem[1016] = 144'h030c0042ff7716adec10f4e61a20e968ef8c;
mem[1017] = 144'he3d11ae8020beb500a791b26e111f373e404;
mem[1018] = 144'h091ce3c0e5b9f4391cbee512eb7101fe18c5;
mem[1019] = 144'h096fe4e61b3c0ac919a5ea9510060f340d1d;
mem[1020] = 144'h17b0f244f5f9f99ef7d2e37619591c131cfb;
mem[1021] = 144'hf7700a6a07521757e818027514ffe697ec67;
mem[1022] = 144'h02321a8d03361efff5410137fefce1c513d9;
mem[1023] = 144'hf386104ced7cf8651dc8e73a0f7004741fd5;
mem[1024] = 144'heaf8f1b9fb26fec8f2551958ecb5f99d08af;
mem[1025] = 144'hf402e2f5e711f8721b28f2581bd7e57818de;
mem[1026] = 144'he2ebf6950af9e485050b182600741ffd17cf;
mem[1027] = 144'hfffa15a9e27f18dff6d60f0d0be706ede484;
mem[1028] = 144'hecd6fc330711052af2afe8a6077b0a0a1794;
mem[1029] = 144'h071ae59d1d38ffa3e899e9ccf45b196d07c5;
mem[1030] = 144'h0fd8ec0af4151fa216ee1fa1f37ffee8e56d;
mem[1031] = 144'hf30bf583155213eff02a12c81b9c1eb00178;
mem[1032] = 144'h0077e8d5fc7ce585f818fd0e0036eee1f65a;
mem[1033] = 144'hfde3f7b0070d047af3f2f0b11a580a29ed28;
mem[1034] = 144'hf552f3c9e4af170cfaf5188e065502ab095c;
mem[1035] = 144'hf6e6edeaeb8006491d0fe6aae89214a9f6fd;
mem[1036] = 144'he04fec9f0a211ffff1111141ee66e09817c5;
mem[1037] = 144'he7cb086b1c03fceff82c1203f63808360613;
mem[1038] = 144'h1257f2dff8c3e62e188de12fe402fba80a63;
mem[1039] = 144'hf74901311b891d2ff0f8105513faf2520862;
mem[1040] = 144'h1fa918fffb85fbf8f71c02e5ee08e567f2fe;
mem[1041] = 144'hffd8edc70bd81e6c1021eee3e8d40980e154;
mem[1042] = 144'h09f3f99bebe5e3d61226eda6ebdee842ed3a;
mem[1043] = 144'h0568084a116afdc01e451ab90cbafdcdfe93;
mem[1044] = 144'h10f21200e5b2f527eda41c11ebbd1ca1e6a2;
mem[1045] = 144'h1397edc7199c1274000a09a9e8090e6f0186;
mem[1046] = 144'h0ab811d316bd00c8149100a2ee65fc5fe1ac;
mem[1047] = 144'hf373f092e791fc31114800abe969e41e0cd8;
mem[1048] = 144'hf33bf9b312981bf204600a96e9360399ea68;
mem[1049] = 144'he2c7ed6a02c8e6c40e0b1006f3c0fa23e490;
mem[1050] = 144'h1efce83112c40123ed1afe0e03b9f108f102;
mem[1051] = 144'he8a70bfdfb00fd6713f31e7be5d4f15ae790;
mem[1052] = 144'h1317fbece4621b8412dcec5c16f0e36cf367;
mem[1053] = 144'hf975fb0904f7f84ffd92f6b60c321c53159f;
mem[1054] = 144'h1ff1fc0fe4830f41eab4e3b1067def040743;
mem[1055] = 144'hfe3f1824e6cd0186f2181965ee40e9a5ff70;
mem[1056] = 144'h049c0136fd62e1c51f111e311ebfe8981234;
mem[1057] = 144'h160201b60550ece609291cc7e2ece6b9032a;
mem[1058] = 144'h11fd0644f28d0a570dbfe752e9b2f2c7e60e;
mem[1059] = 144'h1b2f17640c2b0574e942e1f505c907780f48;
mem[1060] = 144'h076b1f6ff77a0fc70e35fdf115fd15d51263;
mem[1061] = 144'he22d0b6e12baf00b1319ea5608f617a615f1;
mem[1062] = 144'h1ba119df12c1f8b1f55bed23e6f7ea3d0a1c;
mem[1063] = 144'h0254fdc71014fb751a6ee589e145f2030c08;
mem[1064] = 144'h0467067202ee1d490ad3f4bb04670f3b13ca;
mem[1065] = 144'h1dde0685e47c13cae8d1084f1676ff1ae0b6;
mem[1066] = 144'h1e86e143fb18067309ec029c05400576e747;
mem[1067] = 144'h011d172f1202fe41f540e27d13b300c9e7b4;
mem[1068] = 144'hf19efb2bf5230e58ff76053d17e9e4ea14e3;
mem[1069] = 144'h15ae1d60f26f0a641c47ef28e62918140553;
mem[1070] = 144'h1e82ffe212f1fc08ed1de0221f0a1333039a;
mem[1071] = 144'hfebfe0ebfd20118104f9eb640ba61e53e419;
mem[1072] = 144'h1ee6101bfa9f1cfe11ae0e91e18ce32d0ace;
mem[1073] = 144'h015d144d00b20a580f2f09bcf65b08a6ec35;
mem[1074] = 144'h173a1a56e3baf605e919e7f51a09fe85ec07;
mem[1075] = 144'heaa2edd81b58e0bf119614c01d92ecff0ef6;
mem[1076] = 144'h1db7165b1c2812060d1f1bba0dd3e95ef9fb;
mem[1077] = 144'h0796fbb2e5a90798065bf4730c85fa0ce68c;
mem[1078] = 144'hf928041407eb02f309bc087a06ae1b1beaeb;
mem[1079] = 144'he7b104da0e7be950f9bb0afafb23fd781265;
mem[1080] = 144'hf3f717a8fa881c9219ebf79de631eaede464;
mem[1081] = 144'hfbc9ee6ae637f461ffe9f579e44fe689027e;
mem[1082] = 144'h1ca0e8a1ef18ed0d144be76bf658ef061af8;
mem[1083] = 144'hf8a9ec190787e9b3f15c187e12d2e0020b9d;
mem[1084] = 144'he2750ef1fc501c381171eef7e242fa3af0c7;
mem[1085] = 144'h1cb0010fe00cff1ce80308c3f572fa86f7fb;
mem[1086] = 144'hfef00336e0db18a0e8c6fe3fe55c103afa3b;
mem[1087] = 144'h1e6215a0f05fefc20bfcfcfde8c709ae154e;
mem[1088] = 144'hef150327f2ef1aa6fa27e636f93a0464ff3a;
mem[1089] = 144'hfe7a0f611bea0d981aee0feae18bf2ab025d;
mem[1090] = 144'hfdd5f7bc1bf6f5ccf0d20a0507191ea5065d;
mem[1091] = 144'hec6a02dfeeeae7e1e9830d71ea80e213059d;
mem[1092] = 144'h1b2bebfa068bf7d41fd8fa9a0e7f13de12c8;
mem[1093] = 144'he8db0d3c18340b5cec121b760805f65403ff;
mem[1094] = 144'h0146ed73ef28f6f21ddbf3280acaf4230123;
mem[1095] = 144'h0623f26ce926088518e3f4960c2f0146ff8a;
mem[1096] = 144'hf4e20bb50cb00c3102dc09b6133406e2014f;
mem[1097] = 144'h0fb5ec3815de1a0d1abef7cc157000210a3a;
mem[1098] = 144'h03c61e31f71f022b02b4f1281917fa24f2b5;
mem[1099] = 144'h097f1352e336fc221e7f1668e598e22f1cb9;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule