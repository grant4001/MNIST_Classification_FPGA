`timescale 1ns/1ns

module wt_mem2 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h0a49fa2900500251095ffbbbf5770867f69e;
mem[1] = 144'h003201b8f105f7aafada0afd0d1eff6900f8;
mem[2] = 144'hef44f697fa2af612fd54f5e8fd210391fc21;
mem[3] = 144'hf03cf1740610f86af260f32beed0f78cf76f;
mem[4] = 144'h080b0ac1f53e0a35f646fa81f935f83e0c80;
mem[5] = 144'hfb070155041ffc6d09380b7904eb0df5f119;
mem[6] = 144'hf0e4042a0bd00b53f841ffabfc95ffabf03d;
mem[7] = 144'h05b5fd9c060904c30d51f961f670050cf1dd;
mem[8] = 144'hf181f4c70b1f0b77f6bb0a8b012903ef0294;
mem[9] = 144'h0537fe300ad3f0a2f9f7f987f94df57b0848;
mem[10] = 144'hfd0e0935efa10927ffda0d5df2d60bf60456;
mem[11] = 144'h014dfcedef78f1680573f8fdefd0ffa504a7;
mem[12] = 144'hf0ebf7c2f2b30688fda0fd49f3cd08e60ecc;
mem[13] = 144'hf57df8c2f8cbfda7f3e1f46901630ddef0cc;
mem[14] = 144'hf3cb09d10d9504bbf923fd0ff611039d073e;
mem[15] = 144'hfa05f35bef900e21fff5ef46fda1045bff22;
mem[16] = 144'h0e23fc47fe51f7fa06aef82702fa070af620;
mem[17] = 144'hf5ab05acf6fefb8400a1f8490e05f2c0fab7;
mem[18] = 144'hf2cbf8defb210d770b29081a04610513fbab;
mem[19] = 144'hff30064a06b70095f35e091ff18e011bf0ba;
mem[20] = 144'h0aee0a4101fa0c33f0d1fc5302c7f86809c3;
mem[21] = 144'hfab7fc87089b0148f448f910f35dfd7afae5;
mem[22] = 144'h09abfb2ef2fbf17af78c0ba908adf514f8d9;
mem[23] = 144'hf2bc0a8ef9dd076efa4705f6f44afd20f626;
mem[24] = 144'hf414f3cef102f537fd7c09e109d9fa480e49;
mem[25] = 144'hf7c20e8afc9e051d0ae5f5bdf490f3930217;
mem[26] = 144'hfd9a0af10932f5e50ea8f87bf863f263fb58;
mem[27] = 144'hf652efcafeabefb0f98cfacdf11907cb00cc;
mem[28] = 144'h01f6f1dd03460051f4aa008b09cb03c10b2d;
mem[29] = 144'h019bf43defdef9b5fedb05780836f672f373;
mem[30] = 144'h02d3064ef975f11f05a8f79b0eddfaf802bc;
mem[31] = 144'hf4dd0b22f569f0eaf451042ffbcd06ce0a80;
mem[32] = 144'h0a51f982fe7a08fff49306affe57f3600b78;
mem[33] = 144'h0d180c6cfe0104ccfc13044506a0f66bf9c3;
mem[34] = 144'h006ef54e00cbf0e2fa8efedd02db0ef407ed;
mem[35] = 144'h0a95fc14efc70bf4f6ccfe3306c803170f72;
mem[36] = 144'hf97a0e10074fffeff33d0477fadcf28f0321;
mem[37] = 144'h0082f60209e503d60d5e0e8df024f5cff5cb;
mem[38] = 144'h097def8afb4dfa02f9420c0b03390dfa08c0;
mem[39] = 144'hfd48f30cf82a0df0f1d600e2072afdf10698;
mem[40] = 144'h096dfbbb02340450fa550aeff7b5f66605ff;
mem[41] = 144'hf91afe73f704011102f309090b6000eb0747;
mem[42] = 144'hf7f9fad50903057709bbfca9f80201450258;
mem[43] = 144'h08e9f18ef2d1094bfd7f062b03b10b18fb63;
mem[44] = 144'hffbd0a14f4c3ff7af58c065408ad02bd04b4;
mem[45] = 144'hf8b4fd080e03f5940a10094305e8049afb59;
mem[46] = 144'hf42ff0260961fd6bf028f86ef3280c90f2d5;
mem[47] = 144'hf13e0808091b021d04d9fafbffc909f60944;
mem[48] = 144'hfc8defca05970d2d07b3f9f1f0c6fb350942;
mem[49] = 144'h0d3afeb7fde7fb2efb6700f7eedcfff901d5;
mem[50] = 144'h0f41ffd2fa3308e20d0bf425fa7bf5b805a5;
mem[51] = 144'hf3d700ff01c60946fbfd03f40e7f09baffdb;
mem[52] = 144'h0d9af01c0aa4ef55f674069efd46f80a0100;
mem[53] = 144'hf6c70a850b52fc1afd40f16e0f80efbdfb2b;
mem[54] = 144'hf88b00ee0676f678f5820c4f061d00040569;
mem[55] = 144'hf09e0c950a16f9210a7bfd4dfde8f5b3f7b2;
mem[56] = 144'hf330f35a0d74f9ebf5bbfc09f941f86c0c57;
mem[57] = 144'h01d10571fca9fb86021c0a880816081c0d20;
mem[58] = 144'hef7d00f10913031b01e7f4b0f28f03aa02a3;
mem[59] = 144'hf804f7b00811f714faa203d2ff14045c04d2;
mem[60] = 144'h02310e850c36ff16fefcffc9f5dff0d9f13e;
mem[61] = 144'hf8b0fe1e0dfff7080b74f6b30870ffb7f207;
mem[62] = 144'h0917f9320ae3f3fcffc70a0cf9ac0c71f832;
mem[63] = 144'hefb4fa67f02ffabef967068c093003010d24;
mem[64] = 144'h0751ff62f3e5f4f3fef30b3eff6306c60676;
mem[65] = 144'h0aeafe470cd6eece090803d1f6f70a9bf950;
mem[66] = 144'hff62f4a400b3017d06690ce7047907a8054f;
mem[67] = 144'h09e6f3fe0d6cf5d1f1c5ff930721f19bfc70;
mem[68] = 144'h08850be1f525f6370c40f429f3ddf378072f;
mem[69] = 144'h01daf229fcebff7705fc092e0dea046ef90b;
mem[70] = 144'hf547fc72002509790b2af0300b62f56ff71e;
mem[71] = 144'hf2860b26008b0b19010dfa8a0e57050a01b5;
mem[72] = 144'hf745fe1808c7fcc6f271078900a70cbcf54a;
mem[73] = 144'h0d5bffe0fc75f54bf1ccf91e035708b3f1bf;
mem[74] = 144'hf184f124ff80fc440f55ffcbffd2fab8fc77;
mem[75] = 144'h0d8cfa77033809cd07d20ada0fa6f0850503;
mem[76] = 144'hf9ed083af6eef506efad01690558080af1c3;
mem[77] = 144'hef8f0ab9017d01f9025e0796f611f4f3016c;
mem[78] = 144'h0633f062f5b706d7f50201b202a10ab0efa7;
mem[79] = 144'h0a2a0ff303f408f80423fd96f7450fb0fc72;
mem[80] = 144'h0ead0b6f0343f00bf19efa8a0c4fff32f564;
mem[81] = 144'h0397fee1f9cbf0d508dff4ef0425f68ff435;
mem[82] = 144'h0bb0f3ca06330dbdfb3f0a11f13b0ee3fc83;
mem[83] = 144'h04cdf1ec099405cfefbb025af14dfd4cf30e;
mem[84] = 144'hf7fb0d6bf219fba301a1f0f406010bb1f9ea;
mem[85] = 144'hf822f4710ac302b50787f5d8060004adefa0;
mem[86] = 144'hf316ff28f9fbfb5ffd79f4340098f9c40376;
mem[87] = 144'hf5d9fb6403a4f81506dcff85f1630220f85f;
mem[88] = 144'hf0e9fbc0f9b0f689f372092dfeddfbb3f85b;
mem[89] = 144'hf0c3f59d028ef000fe74067f07f4fb6afa74;
mem[90] = 144'h075c0238083d05b1f671fddcf060fc2300c4;
mem[91] = 144'hfc1a086cf561f2a60b27f36c053d08ba0d51;
mem[92] = 144'h07d50255f67e05a809fbf3640cabfe96feb5;
mem[93] = 144'h003b0ba5fa160cc3f239079ef2d2f73b07a1;
mem[94] = 144'hf590f706f330f1d2f5330bc705100007ffc7;
mem[95] = 144'hf95204fd0604f06efacb0db6f4e9ff5df357;
mem[96] = 144'h0886f15cf8ca0d450842f945021ffe280565;
mem[97] = 144'hf033fa59f58704abffeb0f9809180056fbf2;
mem[98] = 144'hf3790796f2a5f2290fa4f8edf7d4f16b0341;
mem[99] = 144'h07520575f2f608bb0ada0a97f695f2f3f6f7;
mem[100] = 144'hf32e082ef770035eff1bfc34ffaf070409b5;
mem[101] = 144'h0013f36b06b3021bf1b3fc91f6b3f0da004f;
mem[102] = 144'h084c0e75073ffcb2053d0e620643f8ebf10f;
mem[103] = 144'hfec0f730f04d0c760e380e4df65bf977f622;
mem[104] = 144'h0935000e069a020a0c2608fcf01802f5f53f;
mem[105] = 144'h0ea8faa7fd87fb0e074208b2fd69f324f94e;
mem[106] = 144'hfd39f25904daf9c4038ff726f6ef0a8afed0;
mem[107] = 144'h0e44fee3f39cff64f90af180ff5c0853f625;
mem[108] = 144'hf49ff8f7049a0b44f5710e73ffd5fbdc0d97;
mem[109] = 144'h067cf6f8f3e101740f6006eb00600df90935;
mem[110] = 144'h025d0c0f071c05d90f1002900dc10ab70216;
mem[111] = 144'h077df1defb81f10df69ff4840ef4f989fa65;
mem[112] = 144'h078afdcaf1ce0db2094ffdd3f1cd0639fd58;
mem[113] = 144'h0a6c0c1401210842fbc9f7cf04b806d9f95a;
mem[114] = 144'h022cf7f404fef77af046fe1409edf2bf0990;
mem[115] = 144'h08f70d54f952f9a3efabf6c0fc610549f056;
mem[116] = 144'hfd5af74bf885ffd90610031d02f00e410b18;
mem[117] = 144'h0c6606edfcba00580ce9f6cdffc9f898f9db;
mem[118] = 144'hff7e0527f27bfe2b0f5e0e8d031a0ac30fc7;
mem[119] = 144'h0a7103b8f36d039000490dbafd60ff4e07c1;
mem[120] = 144'h05fb0757f4eefe68f32df4f00cd0024df477;
mem[121] = 144'h0924f4e3017efa5907acf2c5fc5605260759;
mem[122] = 144'h054c022dfb27f2a7f41f06fcfaca0355f818;
mem[123] = 144'hfc76035cfd88fe3fefe3f29b08efefff055a;
mem[124] = 144'h08c70d54ff8b0525f3690596f1890d6c01f1;
mem[125] = 144'h03d7046d011eefecffd90441027f0ecdfa1a;
mem[126] = 144'h07cef0920003f593fe9a0901fae00a710255;
mem[127] = 144'h0acb0fd2f4ea0ee6066005a404bb0c790154;
mem[128] = 144'hfe2cfe09fd3803bdfccc062f08aff582fd1d;
mem[129] = 144'h05a30d86fea00172009808210963f6fcf8f6;
mem[130] = 144'hfaef021a0a53f24cf5f5027405bdf02cf7c6;
mem[131] = 144'h06c3f3f0f25df97f0daaf1760597fd2dfc9c;
mem[132] = 144'h0d0a032805f2f032f8bd022805a80bbcf4dd;
mem[133] = 144'hffa5066ff2d909a305700b5106abf184fe8e;
mem[134] = 144'h0f44f12bf7a50a12f38c0825fc570fdcf818;
mem[135] = 144'h0d420d6a0c3af56d06f9f5150e5208e2f085;
mem[136] = 144'h04750e61fbd00b420759f4b804c70226fe05;
mem[137] = 144'h06d908f5f54407cd0791f0230399f2dcf7e6;
mem[138] = 144'h06b0f9c404ccf506f7850efa0b28f4480b94;
mem[139] = 144'hfeeb03b3f7070e6e00eef322fe7f0f09f175;
mem[140] = 144'h07bbf2590c36f2a4f06b00e4ff4bfafd0595;
mem[141] = 144'h0f8afe13f3ee05a3fbd60bcb02f0f4f3ffd2;
mem[142] = 144'hffd6f50ff420f07ff21c023df125f0e4f700;
mem[143] = 144'hfb24f80a0cc2f39e079905f107edf3f00bb5;
mem[144] = 144'hf911fbe4fa44fc2cf988fc78017c0edb0e8f;
mem[145] = 144'h08700bd9f469fa4ef2c70504f949f24201d0;
mem[146] = 144'h0c910811f9110b0c0616f8b2f6dcf828fb95;
mem[147] = 144'hf91affd108fa0dd8025efd7ffb56f666f4a6;
mem[148] = 144'h08cb0f60f1f60497fb86f7fcfad306090f5a;
mem[149] = 144'hfe600b2f0b00f0e2f0d1f00b0d54f3120d4e;
mem[150] = 144'hf6e9f85ef8340cef0647070401060aa0098b;
mem[151] = 144'hf514032309d0f0d709eff7f60ef6f16df004;
mem[152] = 144'hfac60adefa6af6f5fd01f9370e20feb50fd1;
mem[153] = 144'h0b93082b0464f32609ee01bdfff70bf90c98;
mem[154] = 144'h0d6bf0a30e87024df9c50b34fe3c09dafc64;
mem[155] = 144'hfd2805110e94feab0d0af20c0127fe2dfa49;
mem[156] = 144'hfbf4fefdfdcbf8e10ccd0186fd55f866f565;
mem[157] = 144'hfe77f0eb0b10fe2dfcdaf5cef822f5bffb37;
mem[158] = 144'hf65201abf682f1d40855fcf7fc71f67ff473;
mem[159] = 144'h0baa00730d13fd630c2e020a030ef96c07b4;
mem[160] = 144'h0126f8710e0cfb35ff0e0ca90358f81700fb;
mem[161] = 144'hf0c5f981f0adfb5705e00246042bf1e1fea5;
mem[162] = 144'hfb9a0c4407e00aca02fd0060f76a05950b36;
mem[163] = 144'hf2a90677066a0367f70d05f1029dfea00cf3;
mem[164] = 144'hfafc014004e8059002e3079f0a9affe30e24;
mem[165] = 144'h01410b3d0d75f4b1fdcff2ddf8f80581fcc1;
mem[166] = 144'h0f5b0b67f6e10a9a008d02a1fa7cf656f93a;
mem[167] = 144'h0516f2370310f47dfea30d650bc3051a0ee3;
mem[168] = 144'h037c00b004e2035f0588f481f8ca0c32f512;
mem[169] = 144'h05a90ed703cef9160ac2f56601c007100b5e;
mem[170] = 144'h06060a920241096a086702db0ab5fe2ff844;
mem[171] = 144'h0d770d420c4f0e72f5bdfad30c06f1050123;
mem[172] = 144'hf63ff92afefbf79c04d4005bf3a9fa2ff00a;
mem[173] = 144'hf6710c16f80303abf370036dfa2ff41e05ae;
mem[174] = 144'h0f3df056fc3ef3df0e360a1efd1b03840a36;
mem[175] = 144'hf73bf8ab042301b0fe6308c20d6803c30662;
mem[176] = 144'h0b3df7bc075bfd76fc6206740702f04bf50d;
mem[177] = 144'hf09906f106370c6a01d80c1bfafbf497f998;
mem[178] = 144'h0f75f4bef544f79d0536fe6defe7ff0d0c88;
mem[179] = 144'hf7dffa9508cb0b8e0dd70950f5290087fb68;
mem[180] = 144'hff4af3cbf9a009020589f7d2f9a0056cfbcb;
mem[181] = 144'hf1dcfd4804b5ff8909dcfc8c05f3097e0bdb;
mem[182] = 144'hfd0706a7f738fe810948fa93ef5c040efb26;
mem[183] = 144'hf3c509f4f37c0b710e22fe81f90af795f0df;
mem[184] = 144'hf730f201f7e4fd7b07ec04bf0e840507004a;
mem[185] = 144'hf8ad0359f334fa780faaf093f67b0753f08f;
mem[186] = 144'h0a770311f541fabff2e4020bf0a900c8fc70;
mem[187] = 144'hfefbf8eb0ee702ea0ec6f195f52cfa39035a;
mem[188] = 144'h0505f76cffc0fde602be0d51fb390841020b;
mem[189] = 144'hff810d8c03e6090702b2f2f608ebf24cfbd9;
mem[190] = 144'hf429f1a6027ff374f2ecf46af347f132fcee;
mem[191] = 144'hf80bf7bc095d047c08630868fbe0ff42faba;
mem[192] = 144'hf76dfb18f6ee062efb5ff120fd84028cfdf7;
mem[193] = 144'h0e0d06270e77f7e9f66e0942fbcb074508b5;
mem[194] = 144'h0e0d0d5ffe3af00a0f50f8c70c270af50552;
mem[195] = 144'h0631f0d10b9802620293092d0c0ef4780b36;
mem[196] = 144'hf305fdb8fb6c0a6df9ef0685f3a00632f7bc;
mem[197] = 144'h01820840fcb0f6fc0919fde502f5f700f1eb;
mem[198] = 144'hfbfa069305e00aed0beef4d60b430f61fbef;
mem[199] = 144'h08ac080f01cdefda044cf8c7f8a40b27046b;
mem[200] = 144'hfb7204ceffc50d5ef8eb09def5d10bd00d73;
mem[201] = 144'hfd10f84900040db2f1cafd500b2b0d2afe2d;
mem[202] = 144'hf45a02a4f17300fcf9860721002a08ed0490;
mem[203] = 144'h0d06f8d4faa9046bfef4f5c7fd34023f0028;
mem[204] = 144'h0610f649f6c301ecf9aa0ea4f5d1f5280eae;
mem[205] = 144'hf8e6f6b4f060fcc107a503520c2a01a7fb1c;
mem[206] = 144'h0d4f0203f264080cf6affe960ceb06b9f188;
mem[207] = 144'h0baf026c069ffadef0b10c0106e40eff09d4;
mem[208] = 144'h059b0412f07efcc5f3cc0c2d0b5afb650f71;
mem[209] = 144'h0084f1cd048afe4bf9aa034901c4040e0d58;
mem[210] = 144'hf7bff80cf9cc012bfc460f6af9900c80f178;
mem[211] = 144'hfa5df090fc27f596fb64f6e004fd05680bc9;
mem[212] = 144'hf08c0b1009630a10ff05041bf045f6680781;
mem[213] = 144'h0ee7072601f6035af5e7f0f7ff64047a0f47;
mem[214] = 144'h0c4bf257fc31f304f34cfbf00eaff408ff80;
mem[215] = 144'h08680245fcedf0640b270ae002370193fb8b;
mem[216] = 144'hf6f4f8e7f693f681fd2b00b9f397f1cb045a;
mem[217] = 144'hf9cbf2210eccf2d8f4c40d9a0d05f1f50cf8;
mem[218] = 144'hfeccf1070e5d00370a3ef0f8058b098e0b70;
mem[219] = 144'hf3d606d9f0c10a2c08f5f58df0850a53fc2e;
mem[220] = 144'hf8290d18fb5d0526f6bf0901fc01fa600489;
mem[221] = 144'hf44a09d30e1407dcf97700810085fc85f31f;
mem[222] = 144'h0c280b9503090c1706e5f574f47109ae0fc6;
mem[223] = 144'h0ca6f79e0d26f462f4dff2610b1c02930ac1;
mem[224] = 144'h06a40ae0f0a3f25d0f2a09cdf92afbd9f28a;
mem[225] = 144'h07dafc70059af5de06c5fe18f65dfe550cb5;
mem[226] = 144'h03a6fb90fef709c503d10f53f578fef20d42;
mem[227] = 144'h05b4ffa0096a05bd092b0040f191f5f2f752;
mem[228] = 144'h0c2b09d1f3cd02edfd96fcf1f55bf02cf450;
mem[229] = 144'hff19fe0cf4cef91cfdc2f6be09070d1ef5a2;
mem[230] = 144'hfe90fc34f218fb7af3020192060c03c40577;
mem[231] = 144'hf2f1f8050d28f512fdba03f1f25f02f6f3e3;
mem[232] = 144'h07fcf5b4efed030efb93f253f51bfaa809fc;
mem[233] = 144'hf4e9041c07cc07d0f0510d710925056bf75a;
mem[234] = 144'hf8bd053ef79b0353031409100a77041af5ef;
mem[235] = 144'hf4cf03e00a7f03a9f849f193f9c0fcd60ebc;
mem[236] = 144'hf903000f06e6f7d6f6a705bc0a0f0561f03c;
mem[237] = 144'hf5c301d40ae004bff083feebfb15f5dc054b;
mem[238] = 144'h0365f4470b4e011d066a03e3fe7207760d5f;
mem[239] = 144'h09dc0e8afd93f8d30d6f0a4d07d900450ef2;
mem[240] = 144'hfb9709ddf777f2c50d3e088aff73006bf632;
mem[241] = 144'hfa38f6e3f030fcd0fceeef500d25fc5c0764;
mem[242] = 144'h016303770e76059b0e75f48e070106eafdfe;
mem[243] = 144'hfbcdfc0e010209d7f9a8fd77f0ef0463ffec;
mem[244] = 144'hfac3f837f2030542f8530e40f9c502e7fe7c;
mem[245] = 144'h096cff0cfda9fd5503cc08110e4b015df727;
mem[246] = 144'hf578fdd208abf3b7f030062806bfff9df66a;
mem[247] = 144'hfab60ee4f45d05850ec80083fbd7f355fbb2;
mem[248] = 144'hf8a10fbb0c290cd30d74077dfb8407ebfc24;
mem[249] = 144'hfa6dfbde091b0b5707d7f134fc1cf01ef8ee;
mem[250] = 144'h054c04e3fbc1f0cdf7dc086cf4e20a97f8d3;
mem[251] = 144'h04d0061901560bfa010a00e901c1fcb301c0;
mem[252] = 144'h0aacfbe5f266f6d40bad01f1f600077900ba;
mem[253] = 144'h0588f32df0c6fc3cfb05f5f40c2a0ecef7ec;
mem[254] = 144'hf070067c01ec0a83f7f8f4acfcadf493031b;
mem[255] = 144'h0bd2f865085cf82df868f962f5860797fcf4;
mem[256] = 144'hf034f34602fc09c1f63309330b050710f615;
mem[257] = 144'hf434fe710b29f7b70819f25900570a9207e1;
mem[258] = 144'h0812f169f82efa070cbe03cdf0f8f03ff4e4;
mem[259] = 144'hf48af034ff0ff69ff93a041df6c5ef3205df;
mem[260] = 144'h055300a0054c01f3025bfcc2020afe0d0f53;
mem[261] = 144'h0e4ef93e0be6f79d079bfdfd01b408c0fbc5;
mem[262] = 144'h02c906eff5630822f8f908a10d90fead0df4;
mem[263] = 144'hf4f306080863ff9909900be4f6ecfd8cfd9e;
mem[264] = 144'h0a260bd0f0fd0a1d0406038df08ceffe00a5;
mem[265] = 144'hf8120f36029f0804f749f479ff4e08680b9d;
mem[266] = 144'hfbfef47df1990b5b09de0c90f355f20c0f24;
mem[267] = 144'h0425f680051b0cb8f9700448fe36f67209e2;
mem[268] = 144'hfba60f2c08bfffa9fd9703e9fa19f99cf1bd;
mem[269] = 144'h004b03a4099bf368ef8ef1a8fbbc0e01fe0a;
mem[270] = 144'hfe950ad1ef9c0cec0a0e0dfb0b250785007b;
mem[271] = 144'h05a4fd5d080ff05a0ef6f4d60001076d0af4;
mem[272] = 144'hfa03f67ef456f05e0cd3fd8df9c30d2e024c;
mem[273] = 144'hf1c6fda1f215f0aafe4ef688f3d50c3004a0;
mem[274] = 144'hff6a072efd4ef6aa05abf3abff27fb49f0fb;
mem[275] = 144'hfa3c0caaf6310154ff5f0c4df811f7aef3c2;
mem[276] = 144'h0681f049f12f0d2afeef0ab5f5930ef9fc52;
mem[277] = 144'h062b089ff9de0e7f0e0bf801ff19fea3f4a4;
mem[278] = 144'hfe7907fef01d0334f15003330836f91cfb97;
mem[279] = 144'h0d16052ffeec0ed5fe5e095dfef9fe3d05a1;
mem[280] = 144'h02cdfd6207f90b54ff320295f9a80b53f7a9;
mem[281] = 144'h01acfe06f6a704a5ff49fec30914085e0346;
mem[282] = 144'hf34805d40133f1c0fa9cfc8f06f8f64bfbe0;
mem[283] = 144'hf545fd790beef649fdadf99df7c50846fab8;
mem[284] = 144'hfda40ad302bf09e5fb8c04a9fd83effc027c;
mem[285] = 144'hf245f4fdef7df1fa0c6607c60f5efb4ff6da;
mem[286] = 144'hf73004290725045ff3f0f16400edf1d0fbfb;
mem[287] = 144'h0cb5095ef1250601fe6effaefca9f428f8e4;
mem[288] = 144'h082cff1406d605d1f87a06de05d50efa0b74;
mem[289] = 144'h0870f066fab30401f322034bfcd00d8d0777;
mem[290] = 144'h08110668f6a204cd07750843f911f07bef67;
mem[291] = 144'h05d1fe58ff2dfcdd00b30edbfa03f0990db5;
mem[292] = 144'h053d0a75fa1f09d9f2960bddf5d608120627;
mem[293] = 144'hef610bf6fe6101d10843f937029ef5dbf104;
mem[294] = 144'hf53603caffd80d35f45ffea9070804a30806;
mem[295] = 144'hf5e805fefb5ff5f50433091b027706fbf133;
mem[296] = 144'hfb79f24af42bf4c806c8075efdb20803f640;
mem[297] = 144'h08e5ff58f241068d048f0d1ef7c00e000c1d;
mem[298] = 144'hfb3b0b010c22f6adfba1f5110ceefcca0f46;
mem[299] = 144'hf371fa70055a0b39f7b30a92fd77f12703f7;
mem[300] = 144'h08d8fe3ffeeef6bd07eb030e0e33f8f2fd33;
mem[301] = 144'h0b77f57af1710b34076502bafd64fcfd0bdb;
mem[302] = 144'h0eac0954ff740398f1320a3af7fbf5f60b11;
mem[303] = 144'h03b00257f20304d70e1a03e8f6dff8950db4;
mem[304] = 144'h0e050eca030ff1bb0419098a0c62f6fc02a0;
mem[305] = 144'hf5d9f08d0f640b3aeffcf3380d930d590c4b;
mem[306] = 144'h0039ffc8fc25f2c906cc071a0e4806930a59;
mem[307] = 144'hf2740ae3046b000304a600cefafaf9e00ac8;
mem[308] = 144'hf4770b030f320bd00ee8f5a1f87dfe41fdc6;
mem[309] = 144'hf7940dc4079807ec02b40692f4d1f67505bc;
mem[310] = 144'h025df6430cdc0b1df40e07e1f94b08590730;
mem[311] = 144'hf8a30cf60ae407810ea2f76e0c9c093df228;
mem[312] = 144'h020a0b3403410b3d0bd0f7ff0512faa70d31;
mem[313] = 144'hf6e604faf90004aaf0930201f375f811f10b;
mem[314] = 144'hf462f708f2f000e90dabf02f0b4809be0ae6;
mem[315] = 144'h028cf277f2a80b99f3740914f9350768f72a;
mem[316] = 144'hf83d0b29f679f9970938035cfaf9f9ca08c6;
mem[317] = 144'h038c047ff8faf2e80ba2032af786f2fc0984;
mem[318] = 144'h0683f48ff52e0765042befa0f93806c8f3a3;
mem[319] = 144'hf770f896f4e1f096f4790fd50ed9097403d5;
mem[320] = 144'hfce1efbdf8df0136ff54f6f60c4df511fb80;
mem[321] = 144'h0de3f3f3f762f0f70f680afcf56bf7230e1f;
mem[322] = 144'hfbb4f804f823fc13fe2e0514049a024ff0b8;
mem[323] = 144'hf27cfa5a070001ed052ef36f0e5d06200d3b;
mem[324] = 144'hf673f55001ba02c0048efdfefad9f4ac043a;
mem[325] = 144'hf6fbffb3f3e9060ef874fd82090200de0a79;
mem[326] = 144'h0bcdf0660681f4eb03510e1efadf033bf920;
mem[327] = 144'hf129ff2d01ea074904970c1cf708f2d7f197;
mem[328] = 144'hf5d60d99f82cf84a0f46fcb7f4b1f6700b3b;
mem[329] = 144'h083cf66ffa77f215f1c6f41b0878f114fe5d;
mem[330] = 144'hffdbff9a0016fda9f96c032303e70a0004cc;
mem[331] = 144'h0c4205a80ecf0adf094df2dcfa03074bf5f9;
mem[332] = 144'hfe5b06ce096ef1490b24f45a0af60007f097;
mem[333] = 144'hfd01095df90dfccffba705e5f1e50bf808b1;
mem[334] = 144'h0e10fd1e101af76ffb6909d3ef04f2e70a5c;
mem[335] = 144'h0dc0fb50005dfa5bf348f41602a70a000ece;
mem[336] = 144'h0e74076ef713fd4b0e4d002cef95fa05f417;
mem[337] = 144'h04b9fdddf74b08a7fa6cf26cf9650702f9e8;
mem[338] = 144'h03c2fa4d0912fd50f9ae05b7f097f16bf6f1;
mem[339] = 144'h0708f8870b9400e502f3f7e508b90946fd56;
mem[340] = 144'hf5e2f6cd08e50dfa01b9f1effdccf6ab03ad;
mem[341] = 144'h0c2c08cd08c608f0fd4008aaf73a03defe16;
mem[342] = 144'hfae8f0b20e7100350b0bfdbbf6b801d903bb;
mem[343] = 144'h0978fd1ff45df6dffdc5f6d9f1c7f0ff0a89;
mem[344] = 144'hff45f41afd95f6aa0391f5dbfec3f79302c3;
mem[345] = 144'hfe1bfceeefd4f022f924f28e0543f100058b;
mem[346] = 144'h012103dc0c8df13efdce00ba0702f8c3f676;
mem[347] = 144'h066cf6e00b1009d30566fbba0a43f9f7fa92;
mem[348] = 144'h0214fd880b4800e600f401fafbe9082ff689;
mem[349] = 144'h0811f4fff255fd0d0516fb9cfd12098b0b26;
mem[350] = 144'hf22409a40b5afd0bf00106860e93071bff2d;
mem[351] = 144'hff1f0f2afdc1002af1de099efdf00b280d44;
mem[352] = 144'hfd590c140d3ffecdfd620985ff1904f709d8;
mem[353] = 144'hfaf6f3fbf17eff340574004e0f8ff693042c;
mem[354] = 144'h0253079e036306ddfe040a3cf441fea7f7c3;
mem[355] = 144'h0d8bf271fe2c025a0d29fd69fa440858f856;
mem[356] = 144'h0d66f6850aedfbeef08c03200836feb6fccf;
mem[357] = 144'hfb70f81d0b3f046f0b0ef0c7f1ba03affa53;
mem[358] = 144'h048104ad05db05e9f47dfce20221f64afd08;
mem[359] = 144'h097af4f3f99f03dc09f5f4940860feb506bf;
mem[360] = 144'hf748fffaf1490b17ff87099ffd3afb81ff93;
mem[361] = 144'hfc3802ebfb02fd78062ff0b4f5bf044bfbb8;
mem[362] = 144'h0ed90909f68a0d62fc0a065cf65affa70efa;
mem[363] = 144'h0970f81ef99403270188f18df9ef0e0efb57;
mem[364] = 144'hfcd50d490627f6b00ab401fb04830784073d;
mem[365] = 144'h0addf85c0a04084bffd703ad0448043d09b2;
mem[366] = 144'h03caf8e60bbcf7bf0c790af60109f13afb8b;
mem[367] = 144'h0717f190fd5406a006b00dd2fe7bf478f011;
mem[368] = 144'hff710a9cf4d50177f040f998fbfc04750e1c;
mem[369] = 144'h06810054eef8009afe67f2110089fc9df30b;
mem[370] = 144'hf929f9de0bc4051ffdf9f9e4f0e9064df1f3;
mem[371] = 144'h0e9205fd09b0fcc60a40086a0dd90e91053d;
mem[372] = 144'hf93ef58604f9fe65f8fc020f0b17007c0031;
mem[373] = 144'h063f03350d3bfc56f4820bb60adf0919f30c;
mem[374] = 144'hf827feadff2907fb0c5c01b80527f436027f;
mem[375] = 144'h0d79060003a3f4e3f05e002e01dbf64afa76;
mem[376] = 144'h0429ff96040af4fcf4aa02ecf8b10832f087;
mem[377] = 144'h029505e001360f440458f74d0fa9f5c2061e;
mem[378] = 144'hf362f93dfcddfc61f946f0a7f7b5fc5203db;
mem[379] = 144'h070f082f01660e8ef54bf55f032e00e4044e;
mem[380] = 144'h0a130e67fd9403def50aefa7f31f02df0a7c;
mem[381] = 144'hf2aaf89b0c650d56ff96f45e0a48f7b7f727;
mem[382] = 144'h0c82f3eaf1350cec08bbfbabfed504adfadb;
mem[383] = 144'h0de8f2250f76ffa00e9f0788fb3ff142f36b;
mem[384] = 144'h030cf440f388f7efff6505edf3240a4e0a83;
mem[385] = 144'hfc8bf62a050804310f4e075b07070126fea3;
mem[386] = 144'hf80bf622f18400fc05a207a7f52d0c0ef1f4;
mem[387] = 144'h07dbf4d9f9a60f4bf183065bfbfd0f37f00f;
mem[388] = 144'h08bdf4b906e40d8a0e9a0cdc04fe01b7fc5a;
mem[389] = 144'h0116f212fdecfaaffd2cff7ffd96f380f732;
mem[390] = 144'h0d3904e403e00dc9f7c208fc0a66f896f08d;
mem[391] = 144'h03a7f8160769f1c6fb2b092c057508640447;
mem[392] = 144'h0598fa7dfa29f7daf21b06230182f52afb2a;
mem[393] = 144'h070007b002490cfa0029f4cefb9dfae3fe8c;
mem[394] = 144'h098d0cfef7820096fec8fafaf64b0ac0f261;
mem[395] = 144'h002e01fff8f7fc29f7070d2e0bacf8f906a9;
mem[396] = 144'h040ffb1e0567f7cdf6f5f2670f8e07820f1e;
mem[397] = 144'hfa41f63f056709adfc550117ffb8fe690409;
mem[398] = 144'h0b63ff17f928fd1afc1d00e1fa7afc0401cf;
mem[399] = 144'h087df96b0be8fb440813085dfb2e0c9bf84e;
mem[400] = 144'h0535079a0136fe2d0189061efc9ffc1b0da3;
mem[401] = 144'hfde605aa0b6c08a4098507f9f58c0b3bfc40;
mem[402] = 144'h0fd3f8d5f3c208e5f7e108970447f4eefb3f;
mem[403] = 144'h04360fb0071b048d0535067b0853fd7bf943;
mem[404] = 144'hfb18fb61f20cf2adf741f13f001a012d073d;
mem[405] = 144'h0207fcdd0cbff42e0b6ef02600a50489006d;
mem[406] = 144'h06e9f235fa14fa2fff100f020317fa1a0700;
mem[407] = 144'hff730f88f4b20625ff7cf9900716f32f0ac1;
mem[408] = 144'hf0ad06c8f50d003dfd600977f89df489000f;
mem[409] = 144'h0c73f0c60d46f082fd2a0cb4f1affa1907e4;
mem[410] = 144'h0c09effefd3af4ebf0a306d20d0cf9e00440;
mem[411] = 144'hfb3ff064ff9bf224096df3b2f1bbf783fa74;
mem[412] = 144'hfe8c0acf0b190ac000a90e0306d0facff8ea;
mem[413] = 144'h00d7f2a2fd3df5390981f94cf147fbbafa4b;
mem[414] = 144'h0490fabefd180631ff01f8500045f3baffc4;
mem[415] = 144'h04ac0bbbf858041b0cfe0cff02ae0b24f490;
mem[416] = 144'hf6bb0a8dfe06ff16089a01bdf23dfa9af2bd;
mem[417] = 144'hf9fd01de0b3809d2f86d0ac9f39ef2eff02e;
mem[418] = 144'hf2d9f7e8f71d07d3fdb7fa65046b07a3fe7e;
mem[419] = 144'hfeee0f1d0d63fb01060a065d05ddffb6ffef;
mem[420] = 144'h0a58fe830a7004b40820f49ef688fbb208df;
mem[421] = 144'hf7e2f4b5ffe7f20ef52bfb5bf385f6c00d45;
mem[422] = 144'h0001fb30fb4405f9056404acf8f30ef706f2;
mem[423] = 144'h01150be80dfd0c19072ffeb3f79cf5080f30;
mem[424] = 144'h091d0309f3d1fe2cf2eb0dcefebb0814ffed;
mem[425] = 144'h057406aff78e02dc0e550232fefff8e7f5a8;
mem[426] = 144'hf7b4f85cf3d800a50df7f01b07d3f249f77c;
mem[427] = 144'hf10df081fb8902c1f9c60bb6020ffeca0f73;
mem[428] = 144'h0f2508c6f17ef6b704270c95f59004f0f2d3;
mem[429] = 144'hfb87f297f56bf44b0144011d06160d010a48;
mem[430] = 144'hf781fbc6fcdafbd8f9a803c6fefb0eca0482;
mem[431] = 144'h00530f280cbf061bfce105bd0f00f8c8f030;
mem[432] = 144'h08f7f8b3fb19fa980ecc07460d0307260d8a;
mem[433] = 144'h004f0bd4fc9d0bdff3ab0c76f6e3f0fbf8a8;
mem[434] = 144'hf8d5fca50322f15308da040d09240ba0f826;
mem[435] = 144'h0964f7fc003efd14f5630295f3710132086f;
mem[436] = 144'hfeab0d720729f43a098ff4a9061f0723062d;
mem[437] = 144'h00f305dbf07ff011024bfee30f550e0ff5e5;
mem[438] = 144'h0246f0b9fbdcf2cd0505fd3d01a9fda9f3dd;
mem[439] = 144'h0443fbedf9b6f3d30e85f016f5b8f114f761;
mem[440] = 144'hfd100d8308eb0e30f32b0758f24105920499;
mem[441] = 144'hff54f397f8edfaaef7ee0c7307570cc100b5;
mem[442] = 144'hf68f0865ef980854f65408b20bc90c27087a;
mem[443] = 144'h0bd00c0e0f7703570c040e170dd7fadafce4;
mem[444] = 144'hfddc09f10ed10dce051a0df2f036fe45efd3;
mem[445] = 144'h0a06f45600520af2fbeafb6408bd00f10bb1;
mem[446] = 144'h0aa706180d22f49c02e8fd9af108fb3ef366;
mem[447] = 144'hf324fbc7f0fcf296f1ab0becf0c4f61c0885;
mem[448] = 144'h061d0875ffd409640a1f024af92bf9fbf849;
mem[449] = 144'h0595039cfa050579f22ef44108350b980d68;
mem[450] = 144'h02fa0456f1f40451f812048ff77c02b2fe1f;
mem[451] = 144'hf3e5f5b9f5540213fc0f06520e5f0edef538;
mem[452] = 144'hf969f4c8fd470511f1a401c7fe6e006a08b1;
mem[453] = 144'h0f96035ffcf40447f9b1fd4f0177ff4e0ad5;
mem[454] = 144'h0dab091b00e4f5280ebdf5b4f1c1f17b0117;
mem[455] = 144'h0b91f11d0b56ff29f54c07baf1660cb9f692;
mem[456] = 144'hf4b3fa80f3bef7c70aa70e70fa880a380614;
mem[457] = 144'hfcbbf8dcf9a0f6d3f88f0aac056eff32002c;
mem[458] = 144'hf8abf311fe390db200ea042ef952f0610324;
mem[459] = 144'h08750cc9fc7a0e66fd600a6b0136f38efc3d;
mem[460] = 144'hfa5dfb2df3d9fff0ff8c0de6ff1e0ee2f5f7;
mem[461] = 144'hf3fa053afa02fd25fe1ef1b40922faf0f70a;
mem[462] = 144'h08850367061d0702efd6f4890a5cf17309d5;
mem[463] = 144'hf2c70f45fd15070f049ef3a606850770fac8;
mem[464] = 144'hfd44f111fc36fa65f74d00f8f74cfc4b08f6;
mem[465] = 144'h0c1cf2d60b960db1ff820ddefc10f50a0d02;
mem[466] = 144'heff0fb01f0f504c0f96eeff5efbf0d470c36;
mem[467] = 144'hfc5202e9054907b3fd26f895015d0eb00c67;
mem[468] = 144'h0bc3051005d601f6f8760ade04bf04610ac8;
mem[469] = 144'h077c095b08a40522089efe7cf026f1c00c72;
mem[470] = 144'h099c0c7a09790ef6fdabf8c30452056dfaf9;
mem[471] = 144'h05af09430c8a0a77070ff0c2f5eef746fb17;
mem[472] = 144'hf306f6b60cb306960971080701a6f4c20448;
mem[473] = 144'hfda1039109e2fe7d0657feea07bcfa550921;
mem[474] = 144'h06c4f3020198f6f8073400eefefb0821fa09;
mem[475] = 144'hffb30c690e53ff9000c0fc9f03d3f3350e3f;
mem[476] = 144'hfa1ff0fff012f52cf88e012805d6f53c0eb1;
mem[477] = 144'hfe7ff7d50245f5cff96b0449f8640000f603;
mem[478] = 144'h0588f7f60626f53e0c64ef5d0c09088f0ad6;
mem[479] = 144'h0faafc010ceef6210b91091200cff177f051;
mem[480] = 144'h00def6e2f62703f7fcedfcd50fe902cd044a;
mem[481] = 144'h04b5f8d70e8cf9a4f0830202001f0332fcab;
mem[482] = 144'h0f70ff1ef0d5f6d7f0aefa7ff57f0119f476;
mem[483] = 144'hf227fa20f3c4f82df757097df394089300e4;
mem[484] = 144'h07f3fa4c05e4f858f200f34f0499f2aefa88;
mem[485] = 144'hffa70ce4000c06ee059a08390d0ef3020279;
mem[486] = 144'hf0820ea8fd9d0f0f0c91096b09d209890918;
mem[487] = 144'hf184f352ff970c84073801e9fe75f57ff176;
mem[488] = 144'hf82ef2c80335fd0bf4470c3a05da00010e62;
mem[489] = 144'h08350e89f0bcfdab0be2f74600a9f62706a5;
mem[490] = 144'hfd2ff08a02cd0e1b031c05cffeeaf0390c8f;
mem[491] = 144'h08020d290078ffe301c7f059f3cf06d2f072;
mem[492] = 144'hf1b1049308e1f3af0705f0c90800f1e30893;
mem[493] = 144'h08e9fc4203d40930f7d90290f73803e3f6d1;
mem[494] = 144'h0e01082cf914f912fb16fda0f548084bf059;
mem[495] = 144'h0d86083df8b0f9de0f0607ccf04808d8f5d8;
mem[496] = 144'hf862ff99019c02830c100d7b00da02fef7d8;
mem[497] = 144'hf8dc0e0800b0f8f5f62efa580463f3a10035;
mem[498] = 144'h0cf40a7a039ef7dbf524fa7ffb940b55faf7;
mem[499] = 144'hf245055af8340aaf063f0423f444f92af0fc;
mem[500] = 144'hfd7df3f304d10405f309fb060219f99c0c78;
mem[501] = 144'hf77f0934f2a50567f6c3ffbdfac10518f966;
mem[502] = 144'h022307f202bb0291f43c025afb0f0b940a0f;
mem[503] = 144'hf7b70c51f315f9cdef5ef10df3560c87fae5;
mem[504] = 144'hf7830aa8f4af015d0be1f314035d025303ce;
mem[505] = 144'hfbf6f503085cfdf2ff20fa2ffd73fc7006df;
mem[506] = 144'hf94e0c6203d1efc7019dfc98f9a6f6500357;
mem[507] = 144'hfa500965f50b0a27fe1bf47bf80ef7a0f146;
mem[508] = 144'hfde006530cfb0d88041d0c21065a0e24f92d;
mem[509] = 144'h06a90df2fd7807d0fa73fdfef874f103efa8;
mem[510] = 144'hf7d303c7f964fcbdf39801480df603fcf740;
mem[511] = 144'hf9010d79fcfef55a028effee0e6a048cf408;
mem[512] = 144'h010ff2510ac0f91cfb52fe15f70f036df8a2;
mem[513] = 144'hf268fadc0e010c4f0ae20b2efaf0f93efddc;
mem[514] = 144'h0ef0011ffc20f41cfef4f1abf26bfb2e0171;
mem[515] = 144'hf5f0f96e03b401f409fef485ffc9085ffb62;
mem[516] = 144'h001e065205a1effef1d4fe630c2c0bb0f175;
mem[517] = 144'hf9f5f3e0fae9fcb7efb0fcacff940b2efe59;
mem[518] = 144'h0db30232081e0ba2f32f00f20eacf6450adf;
mem[519] = 144'hf30103bffef7fdbe0310f0820dc9fcdefb67;
mem[520] = 144'hfd76fc360c9ffab3f95d04e0f934f7660985;
mem[521] = 144'hf9c50283f6d8f7e1f5550974faa2068906d0;
mem[522] = 144'h0f820894f1140bc3019c08b30375051f0b55;
mem[523] = 144'h080f0d90fa5af2a2f0e101fbff210e9afa5e;
mem[524] = 144'hf921017ef4cffa47f88bfd5209920acb0ac3;
mem[525] = 144'h0d840bf1fb86fea2fdf1f930032ffa26081c;
mem[526] = 144'h08fafc9ff4270432ffbbf8c4060d00b90875;
mem[527] = 144'h0884001af0180dc50e33fb9efbebfc6bffeb;
mem[528] = 144'h08a403cefb91fa87f27c00bcf8c10a93f18a;
mem[529] = 144'h087c0062fd4c0bdef5460def0deef8c207ce;
mem[530] = 144'hfe38fd5a00790aaff389f875f928f4020b70;
mem[531] = 144'h0a8afdae098703f4f9c6fa5af478038e0c17;
mem[532] = 144'h022a0b21f47efb44f8a3f90701f2febbf015;
mem[533] = 144'hfe3df3c6f09f0387097f063c000ff437f58c;
mem[534] = 144'h016409f1f18cff1bfe850a3a00110e81f1df;
mem[535] = 144'hf8f00b920ef7ff5f092ef791095d00740e06;
mem[536] = 144'hfe3d0bcdfb35f8fbf23201cb0d7cf3fd0b0d;
mem[537] = 144'hffaef6970e3df022f9f80019fa830d2e04f6;
mem[538] = 144'h077bf4ff0946f49cf09401bbf57ef5ae05cf;
mem[539] = 144'h0863f80a0795f520fae30db4ff73fa98f411;
mem[540] = 144'h058bfa1f09c604a40ec1f71c0a5ef1aefee9;
mem[541] = 144'hf24eff770485f2f00caa0022f5ac00cb0e12;
mem[542] = 144'hfc5ef4f7fbedf801f2ec0c21f95eff48f1d5;
mem[543] = 144'h0e3000fb0648fe0cf3bc032f0c890b130b41;
mem[544] = 144'hfe94f465084ef4dc01f807110a70f406f0c8;
mem[545] = 144'hfb0a0e72fc3cefe10f2efed60c75f1fe028b;
mem[546] = 144'hf5cd0448028af9f0fad1f2f0f438fedaf474;
mem[547] = 144'hf57a0613f0f601abf00802a1f723f3720f7d;
mem[548] = 144'hf76df509f96ff8e4fd4d0d58043cfedcf144;
mem[549] = 144'hf558044ef028f6f6f12cf62cff5a0762ff97;
mem[550] = 144'h0354053e0a6af4780665faef01070df704e5;
mem[551] = 144'h053006ab0a3df2c200da0657f4f3f0bbf755;
mem[552] = 144'h0f89f370fa71f8d4f733febb0cc0f904fd05;
mem[553] = 144'h0c03f2480e54fa2b0f6f0cd0fdbafdecf109;
mem[554] = 144'hf81e0fd20a350d950c250e61fa54fc90fbbd;
mem[555] = 144'h08ff092bfbee02de01fc04770fcb0aa0fa9b;
mem[556] = 144'hfe38f055fdedfbe8f24bf1f802b7fd32061f;
mem[557] = 144'h02b6f2cdf45cf343f69601600a18f09d09f7;
mem[558] = 144'hf561f21af6a00aea0c6efe87f8eaf2720071;
mem[559] = 144'hf2fcfafd0c22039dfda9f66a01a90b010094;
mem[560] = 144'h0ab0080af796f11ff007f42bf9d9fe6cffef;
mem[561] = 144'h0de50746f10ff0ff0ae506350ddbfe50033b;
mem[562] = 144'hf0d3098ef209f78c0174f12c0233effbf7db;
mem[563] = 144'hf576ffa5088905fdf490f89906290cb10428;
mem[564] = 144'hf8d4f6c6f49c079d06b3f4830356f4bc00e9;
mem[565] = 144'h0c2209050b65f91301f00ca1069dfe9ffc0a;
mem[566] = 144'h0312f114f870fdb604b4f3910ecdf2f4ff96;
mem[567] = 144'h0b0508c20ac4f06f0dd8f92905d0fd1d0d28;
mem[568] = 144'h0b050229f93906fa0309016efe0a0304095e;
mem[569] = 144'h04cb0820072a03aa06be059402be0172f4a2;
mem[570] = 144'hfefcf53d008ef94c0f100f17f0c90b6ffe9e;
mem[571] = 144'hffc7037df9cdf81af9f1f092f956f865ff2c;
mem[572] = 144'h0c8b0a450c56073afbc1f0b602df04a40951;
mem[573] = 144'h0b330c99fb2802bcf33c044bf90cfc0ff232;
mem[574] = 144'h06abf73af8f2fb4af406040f0011fda3065f;
mem[575] = 144'h05e7f5c2f80b0ed0f46906d3058bf10f0dc6;
mem[576] = 144'hf235f487fc1109fcfdfbfe1002d9fefafc17;
mem[577] = 144'h06530953f5cbf3200b5906d30523efd207ea;
mem[578] = 144'hf16bf61af8b80d710f500901fa71f5c8fd17;
mem[579] = 144'hf3df0945037e072bf706ffab02fdf12c0931;
mem[580] = 144'hf23d0692f374f65f086c0c7d0c1d051afb04;
mem[581] = 144'hf864fa4defc6ffcff1df0be7f64f011f017b;
mem[582] = 144'hf0d4fe610718fcb30a12034ff0d8024dff8e;
mem[583] = 144'hf0f201a9fefffb94fae9fb7df1d201e50255;
mem[584] = 144'hf2410cfb05d2fccffe8efc23ff55f753f91f;
mem[585] = 144'hff2a02c5fe17fe0cf5cb06c6f6ec01820e36;
mem[586] = 144'hf4fa047a00790a760809fcd9f33b0ce80b5a;
mem[587] = 144'h03bcf3dd0fd20d18f4ba0f28f45afac0f372;
mem[588] = 144'h036f00ad0b35ff80fb9108e20b2f0968f680;
mem[589] = 144'hfc82049df546ffdbfcccf07908930628f842;
mem[590] = 144'hf818fc0a0a89f9a403bff08bf680f5e40508;
mem[591] = 144'h08fd0f57fce70ac5faaa0056036c0cdafb09;
mem[592] = 144'hfdd30805f06cf2ed029ef4f2f08709b5f1c2;
mem[593] = 144'h0c260311fa790c9d0d6104d0f54701daf203;
mem[594] = 144'hf30d00930e43f5a70c02f130f0c706e10660;
mem[595] = 144'hf6ba0d7601fb00600447f674fe31f661f128;
mem[596] = 144'h09840d9cfd7e0b71f06df976f44609a3f2d3;
mem[597] = 144'hf4590262fc1cfc9d0e830acb01a5004904c8;
mem[598] = 144'hf1f2f74affe9f7a008fffb660bc70d32fe9e;
mem[599] = 144'hfaaefe85033dfc08fb44fbbe01bbfe96ffb1;
mem[600] = 144'hf0f40c610f7208b6f605fca6f13c06410734;
mem[601] = 144'h0e10f3c906690630082af12c08d90dc6fe21;
mem[602] = 144'h07150b7df03c0e7f09410261fb71faa70489;
mem[603] = 144'hf862f06df46af70ffae6f26cfc00f7280f69;
mem[604] = 144'h036ef375fbd002f7029606540f3bfb2afbaa;
mem[605] = 144'h0ab5fcaf0856f826f7d709c2fe09f326f792;
mem[606] = 144'h02e7078d0f500541fe3ef8b0f9180a9d01e6;
mem[607] = 144'h005af06ffa810886054bf2580d820cdaf16d;
mem[608] = 144'hfb5e0dbe01b9058bf6540abf00b30781f129;
mem[609] = 144'h050f0a57fa700263ef8409b7faee0de5019d;
mem[610] = 144'h043c03500bddff23045f0ed50d83feedf35f;
mem[611] = 144'hf572fe47047e0e30f19c011ffa8ff4ad09cf;
mem[612] = 144'h087bf21807bcf8410eb6faaaefbd0197f83c;
mem[613] = 144'hf80af408f78700a4f9260cb3fd61f24f04c5;
mem[614] = 144'hf6870016f9fa015afa31fa81fcf6f958fee5;
mem[615] = 144'h09bf0803fc70f3eaf553fdfcfa2bf0a7f719;
mem[616] = 144'hfce606610297f3070ba90db0f9ebf65e065c;
mem[617] = 144'hfd7bfb3e04a9ffca06950885fb31048ff5b3;
mem[618] = 144'hf5f4f1bf017509bd03b5f436f47601be0913;
mem[619] = 144'h01e80aa0f3ef03bbf51009190adb01df0384;
mem[620] = 144'h0bceefcaf7a1fd5b0a62fbe50617f96fefdf;
mem[621] = 144'hf6f0f90b00ee0af0ff8dff310a9809960d8a;
mem[622] = 144'hf599f856f6bff126fe21ffffff76fc880411;
mem[623] = 144'h04a8fa38045df1200a41f799f993077e09eb;
mem[624] = 144'h02500ce40774ef7dfdc9f60ff11d012e0f72;
mem[625] = 144'h081bf830f1490b120926fad2fcecef87f60b;
mem[626] = 144'h0ca1f7c2f09a019e0dd1ff35f297069706dc;
mem[627] = 144'h0eddf1baf987080f089ff389f2a2f7e20c84;
mem[628] = 144'hfe6e066ff26905b10c19f0cb0a68fccff73b;
mem[629] = 144'h07f70c88f68ff384f3e3fe640dcdf9a1fd41;
mem[630] = 144'h0eca0671fe7cf7c6efb9ffeaf0a60f5605c7;
mem[631] = 144'h04acf89df9b6f5a8f05d0f00f3a501fefd9c;
mem[632] = 144'h01f2f8f3ff8bfcc80bb9f8bbfc3300e30910;
mem[633] = 144'hfdcf0d820229f8ecf98807320544f5e70533;
mem[634] = 144'hf2f005e9f43c01c40712064ff746009207a9;
mem[635] = 144'hf32afc99056b09f2f1c1f3260c8100e2fadb;
mem[636] = 144'hf352012b025ef98804b300c7fa6ffd20f80a;
mem[637] = 144'hf336f4a60e6a0700faea05f307080e710d21;
mem[638] = 144'h04ec0ee3f927fb21f6a5f161ff58f8e4f535;
mem[639] = 144'hfb88f5b6f03ffde00e61ff53f4d2f5aa02d0;
mem[640] = 144'h0e1bfb030dc809f2f3f403430ad30099f3a9;
mem[641] = 144'h0df1f4c6fd4e0dcef872f79afaf801bcf3bc;
mem[642] = 144'hefe40282fe4cfb8ffb55ff5f0d9afc08fb6b;
mem[643] = 144'hf27af23404f40b320992f374ffeef35d027b;
mem[644] = 144'h0c59fe2ff5fa05f3f8f80b340bf60499f830;
mem[645] = 144'h0993f28cfed0074bf1e4f242f789fe59f856;
mem[646] = 144'hfc400210ef8cf0900f4309bd007e0263f7d4;
mem[647] = 144'hf6df0a3a0d08f98105b007a9f74f0ceb0632;
mem[648] = 144'hfdf3f678067b015af2de05f10fb3f4ea03dd;
mem[649] = 144'h0ee4f67bf7ecfb53fc6cf1b1f1f705f1fdec;
mem[650] = 144'hff3004020670083804a60682f2c00ff10a29;
mem[651] = 144'h0c56068e02b7081a0c01f8cff654ff69ff10;
mem[652] = 144'h0537f3320d9f0d4af003068af6b90ec0f24a;
mem[653] = 144'hfc0c097ff42f0b73043f0dc700a4ef5601c4;
mem[654] = 144'hfdc2fd98f215fdd304ff08cd06da03d906c9;
mem[655] = 144'h03df0dd3faa60195fb6df838fc2f0dddf717;
mem[656] = 144'hf424f7aef0430c950b1e08c7f060f05e0a5e;
mem[657] = 144'hff5b0f3bf87ff0f403c505d8fae909270475;
mem[658] = 144'h00f8f36802d0ff5d0d83fba4fc74f42203af;
mem[659] = 144'hf13406aef2660edaf2cf0e4dffaf0c98021c;
mem[660] = 144'hf786eed90d58fecbf1e6077701aa05fff510;
mem[661] = 144'hf2f6070903ac06800da1f62dfa4afd500875;
mem[662] = 144'hfdee0cc805260c42f413072bf946042301a0;
mem[663] = 144'hfcbafe900ec8fbb003d3007df5e30692ff76;
mem[664] = 144'h0039f3e2f3420834efa500f5ee9affc7fdc9;
mem[665] = 144'h03c3f0dc080def57f876fa2c0df90a14f46c;
mem[666] = 144'h0210fd4cf7f9fdb60d270da909b9fb970b0e;
mem[667] = 144'hfa1ef843fde5f2cef16d02790ea309910bd5;
mem[668] = 144'hfdc20afa017b0e3b0b2807a00946072cfc25;
mem[669] = 144'hef7804010797febf0a5efc04ff340087f610;
mem[670] = 144'hfbcd0c1908ce019e09f80239f678f606fc17;
mem[671] = 144'h09ea003009ea08b4ff08f3c1f816fd9101d9;
mem[672] = 144'hfaa0fa7f049d000ef5a20cde0d34f00707cf;
mem[673] = 144'h059ffad7f8a3fdb3f54a0788f0ab0c3af7ef;
mem[674] = 144'hf7a608b30a54f39b0f3a0f4bf50c00e4ff3c;
mem[675] = 144'h04e603db08350517088befc9fcf0f49a0252;
mem[676] = 144'h0c4d06060380fcf7efcffedff90507c7ffea;
mem[677] = 144'hf58b056cf0aafc04f586f6410cc60b2200b5;
mem[678] = 144'h08c20676f4950b910549f6850f0eefe304d3;
mem[679] = 144'h0a3df102039dfe790549f9b3f44b02bcefb3;
mem[680] = 144'hfb730e590ebcf64ef01c0769054df0d7fd15;
mem[681] = 144'h0780f544f832f24a082a08290238fc85fe53;
mem[682] = 144'hff500a340eec0c67f69f0679f426fc9cf30b;
mem[683] = 144'h0332f3ae0442046c06bb0092f4faff72fb6b;
mem[684] = 144'h0c7f04de0155f4dffb77efadf4edfd960a4f;
mem[685] = 144'hf4e2fce5f675078b0302f4d1039608a5fb39;
mem[686] = 144'h0554f9df0171017b08dbf6e6068bf3d60af9;
mem[687] = 144'hfce0f8dc0b48066ef9ff02b80d150bc6000d;
mem[688] = 144'h0f3d0e12f99ff21ef108f7ec01990f440a77;
mem[689] = 144'hf6b506e1fe4ef02bf74ffa0e04690b6dfcd4;
mem[690] = 144'hf474f33303880ccb0eb7051e08910b160603;
mem[691] = 144'h0a5e0c2af1fcf924063a0fd4f02804710a9e;
mem[692] = 144'h02bcf41208e6f9e306f7f6360a800c65f341;
mem[693] = 144'hfadbfdc0f041f4a6f8d2fe0b007404ecf46f;
mem[694] = 144'hf1c0f5d9f1e3f3dd0b320ab8fc29fa67f1b7;
mem[695] = 144'hfd3e0aca0e1cfa66036208450a4b0edb08d4;
mem[696] = 144'hf9a1f0ccf78804470017fb9101930ea4001f;
mem[697] = 144'hf24e0b7b0d3d089cf303fb95f9aff2890496;
mem[698] = 144'hfcff0ff8f31af57afe680439fc37081900b0;
mem[699] = 144'h092d00fd0e76091c0780f3690fbc0972f3ad;
mem[700] = 144'hffa4f61204c80adfff47fd57fb82fffa0907;
mem[701] = 144'h05bf0718f3080ee8f9a8f49ff68dff96fc4f;
mem[702] = 144'hf9cbf566f65ff5a2fe1df216f065004df002;
mem[703] = 144'hfd1604c10c7b0f9dfc4b0913054dfc82ff5e;
mem[704] = 144'h0c6cf903f8e0f052f525fffd0c9df8ebf173;
mem[705] = 144'h01050f12fc890988f4620bdbfac30b2cfc9f;
mem[706] = 144'h009cf5a7f49df7d30319028ff6b204430522;
mem[707] = 144'hfc2e02a2f79e0ecdf90ef80306f1f43e01e3;
mem[708] = 144'h0d8803b6f7de08eff0cf09b9f3f0f48ef1e8;
mem[709] = 144'h0dff0d8f0df3f104efb4f6c70711083cf174;
mem[710] = 144'h030cfb5ef089fc5104cf094ff7700e7df538;
mem[711] = 144'hfe22f92ff25200f0f292f39e04c4f6540bb2;
mem[712] = 144'h08aa0e7d0ee90f6102190b0101000259fb96;
mem[713] = 144'hfbd806eafd8ff252faa60d0ffe53f0faf3a5;
mem[714] = 144'hfac9fec80793fdd0006f0325f1e30a72f893;
mem[715] = 144'h09dff0adf07afe7907d00d0300090a710268;
mem[716] = 144'hfa70f42f04adf7cafce5fcbbf92407f60118;
mem[717] = 144'hfccf0670f21504a70033f623093efe4dfede;
mem[718] = 144'hfce5f02006c6f26b02dc043909fe00fe0a2d;
mem[719] = 144'hf47bfd630a84f3cffa3601b10b4c04f3f5a7;
mem[720] = 144'h0c36f112f1eeff000a71fdd2f7e4fafefe3c;
mem[721] = 144'h09dd0974f920f107fccd09fd091d0a8f0643;
mem[722] = 144'h0606ff4dfba3066af592f95af92f0927ff30;
mem[723] = 144'h07790d3df216f481f6acfb2404c1002ffa51;
mem[724] = 144'h0530fd1e08ccfe220df403f3f8b0094df30d;
mem[725] = 144'h0c000f5b00f90eb90bda002b0374f00c0ed5;
mem[726] = 144'hf372f516001206bffeabfadff15e03a2fddb;
mem[727] = 144'h0b64071affd4f0dc03ad001b082eff730e33;
mem[728] = 144'h07cff822019008f3fdadf352073dfe590730;
mem[729] = 144'h0c250f7df284f98803e3f547022e0fbaf7b3;
mem[730] = 144'hfa58024ff84307b2f01af177f6f803d20058;
mem[731] = 144'h0fdcf8e9017ff431f239fdd9f577f72f0ad2;
mem[732] = 144'hf058f5a7f9d4f1c8fc430e25088df42009fd;
mem[733] = 144'hf6750ce3f70dfe8006b3f78207bffccbf51d;
mem[734] = 144'hf67601f201500410f5bd06b70f72ff6bf831;
mem[735] = 144'h07c103b30f520ae700f90e360108f5c80194;
mem[736] = 144'hf8b6f0fdf149f4e4f93d0469097008830712;
mem[737] = 144'h096ef1aa0ad3fc26f82d0b5f050b0aa1f438;
mem[738] = 144'h060cffc8f32200aa09920ec40b2ef22500a8;
mem[739] = 144'hf889f86506f90f980bdf0b2afccaf08dfcfe;
mem[740] = 144'h00fb085b08980006f205f54f0a3bf7cb06b0;
mem[741] = 144'h07c4f477f9880cad03cf0a40efd4f630f919;
mem[742] = 144'hf32ef80108840df4fb69fab10b7502a10961;
mem[743] = 144'h0157f65b0f3501c70995f67507abfd69f474;
mem[744] = 144'h03d8fbacf5d905b2f6fff01d026f044b02a1;
mem[745] = 144'hf8e709b5ffbe0351f3bffa6801ee0095fc04;
mem[746] = 144'hf88b03f40b2b0a71f53908c80b9bf777f535;
mem[747] = 144'h050bf475fc86f26d0122099c0b9c0e5afd9c;
mem[748] = 144'h0edef0c7fa05f677fffdefd20d4106460c73;
mem[749] = 144'h0560028f0e9c07d8056c04410beff82c0258;
mem[750] = 144'h0954fad309360acef1610b360ebcf6f3ff1e;
mem[751] = 144'hffc8fca3fb41f5530cea00e10f80070bff92;
mem[752] = 144'hf358f2520b70f3750490f94f0e6f020ef43c;
mem[753] = 144'h0e7e0e54fadff906f8acff98fc1103e004f7;
mem[754] = 144'hf782ee1c03f609d9fb74f7220183083a0551;
mem[755] = 144'hf03cfe4c000407970c4ff8c60f00f4a3faa6;
mem[756] = 144'hfdfef3e701ba0baeff7b0a44f9c1f81204d9;
mem[757] = 144'hf7b5fab9f6c6f429f872ff850cf6f32df432;
mem[758] = 144'hf2fdf3680fd1f0efef46f3db0d3bfa35f019;
mem[759] = 144'hfc62f99c06580e0bfe1df5470664f241f664;
mem[760] = 144'h0de80bf8f4dbf1290972f07cf7f70b5a0351;
mem[761] = 144'hfec70c760a72f6adf04304ae09a4fe7dfa49;
mem[762] = 144'hf1f9efa9012907e20dd8f5d700c804150090;
mem[763] = 144'h0f20012ef10c0f64f696f582f7aef456f089;
mem[764] = 144'h0eacfc4cf10401f10bd00146ef9602ad0b2c;
mem[765] = 144'hfc50f2da03c806e3f89800950a6d085ff87f;
mem[766] = 144'hf92f01b2fb37ff44fabaf5fbf58100c5fe43;
mem[767] = 144'h04f201dcf132068cf01309f80cd80575f7f6;
mem[768] = 144'h067afe2802180f290c9dfbcf0c4a07a70dec;
mem[769] = 144'h0b600adffb63f8d80dfcfc48fc40f240f772;
mem[770] = 144'hf3fbf65307f2fdad09ba0bb4ef27fa4cf266;
mem[771] = 144'hfb8a0941f9a8f50905f300e6f83009c5faed;
mem[772] = 144'hfc6dfd48f2f7fbb5f672f0880a040d3bf714;
mem[773] = 144'hfc0dfa27fbf7f4030bcdfecdffa80d910725;
mem[774] = 144'hfeb106e40b430edef1f30d9e0c89f5fefdc1;
mem[775] = 144'hfa9af5e2039ff4e5fd2cfed607a4f2de0a23;
mem[776] = 144'hf061f103faf5f37bfcc2027804120ecef60e;
mem[777] = 144'h0df80105f7260d7af532fdfe01fdf4c3f590;
mem[778] = 144'h0459f9d3f428f8fff291faea062e0e43f815;
mem[779] = 144'hf33c07b1f790f11f0fcbf223f85309a20f95;
mem[780] = 144'hf79dfb3ff2fef45603240172f4b8f109f5e7;
mem[781] = 144'h049a06b20aae0d54013cf4e50645ffa8f1f6;
mem[782] = 144'hfb1b0677038c0ca7fc55059af2a7f5060ef5;
mem[783] = 144'hfd2a02ce050b045d0ff4097203af09e600e3;
mem[784] = 144'hf0210b990dc70eb50f29ff120f55f220f9a1;
mem[785] = 144'h016f01ef0cf90fb1fa27015f0c90f0230b18;
mem[786] = 144'hfd910d1504100874fb30f92a0eaa00150ccb;
mem[787] = 144'hf31cf4240a470e48034ef12ef0de09e90811;
mem[788] = 144'hf54207f3f69ffa87fd6aff36f88efd5ffe81;
mem[789] = 144'hfcbcfb58f3db051a09680d1a09dc0a42fb87;
mem[790] = 144'h09530178f52ef585f56df8fa04590af9f3f5;
mem[791] = 144'hfe25fd74027504bb058d08ecfce70bee0675;
mem[792] = 144'h02fe07b305ae0cb606d70c8501640b310636;
mem[793] = 144'h06d407e3001cfc7df35cf591069c0656faef;
mem[794] = 144'hf2c2f4a10002fe8408d10a5c00a700be007b;
mem[795] = 144'hfeb304b601500b59f7b8f11202dc00e4fc2b;
mem[796] = 144'hfd97f789046a0d73fa1ff8feff2dfaf70eb7;
mem[797] = 144'h04fd0d06f6dbfa0802d9090dfa450b3ef020;
mem[798] = 144'hf35af8aef5cd0069fcd2fcee0b5ef67e0fbd;
mem[799] = 144'h03c7fe120562046f09780cd9092b09130c19;
mem[800] = 144'h047cf9a109a9078ffc9df8affd0804e2f4e7;
mem[801] = 144'h0131f3e70c70007efa7afa16083afc150cae;
mem[802] = 144'h02f8f18b00e70443f39e069efb6ef4b2f874;
mem[803] = 144'hf52e0e2ffb15ff6709fff0ae0544fa19f7f2;
mem[804] = 144'hfa430c56fa8d083eff310aa90655fbbd0d1b;
mem[805] = 144'hfd9c05f603b20378ff34f21f0ac1f0f70a7a;
mem[806] = 144'h04db011cf5220d58f03af894067ef169f029;
mem[807] = 144'hf62cf5120193fb370cd2f73f03fff9be00e1;
mem[808] = 144'h07e3f8f201cbf803f9dcf53303d4075cf3d1;
mem[809] = 144'hf2a3046af121f94bffeb0d6cff6207220097;
mem[810] = 144'hf676f145f95304ce01c809dbf70af4caf05c;
mem[811] = 144'hf997f5850c07fccdfc1cf33606ae09c00501;
mem[812] = 144'hfa3ef5660bee01f502e2f305f251f8ecfcfb;
mem[813] = 144'h0bf20a030a8ff59a0229f529eff40bb8f403;
mem[814] = 144'h0c66fd4efb4df8d705860a89f0ecf4a4f288;
mem[815] = 144'hfcc3f85c0dac0d650ce80cc30f85f657f746;
mem[816] = 144'h099ff622f733f2e0fed1f579f83d06570e4b;
mem[817] = 144'h0711feb30b5bfb60031701ee0170f5dc02f8;
mem[818] = 144'hf6590c3804580a4a00140ef9fa95fb16f958;
mem[819] = 144'hf13cf28ffc4bf298fc26f94b0eb6f8ee07cf;
mem[820] = 144'h080a092ffbf4020fff2306f902100e7709e8;
mem[821] = 144'h057cfe99fa3df60804eafa710ab2f89703e9;
mem[822] = 144'h0e9c06750d0cf41602cefc52fceafb40f7c8;
mem[823] = 144'h0c4a0e56f0cd04f4f0f304860e70064ef987;
mem[824] = 144'hf67dff60f3aef40ef09f0d84f0620230fab6;
mem[825] = 144'h0da00bb4f949f5c5f0f502edf8bd0f0b09ab;
mem[826] = 144'hf5e3f031f5abf0c2fd340151053d0db0043c;
mem[827] = 144'hf5dc00c1f90401bbf35903cbfe15f3e7f052;
mem[828] = 144'hfd490a5efe60fe03f6baf3bb00f2f8c60c1c;
mem[829] = 144'hf99ffde6fcae07c50c2105bcfd68fe0907b1;
mem[830] = 144'h0dc7fb9501370749f5a70c8100e0078d0b5e;
mem[831] = 144'h084cf732f6e60c78fdf60471030cf133f262;
mem[832] = 144'h04c7fae40b870f3ff8c2f057068b00fe0d55;
mem[833] = 144'h0acd015d0de3ef2af9b8f1610ba6f760fcce;
mem[834] = 144'hffc20506f12804b5017a0e900f080d8c06c2;
mem[835] = 144'hf8700009064201e20f91f8a801230bb8f819;
mem[836] = 144'h01180edafc0af874f72c0bf0f60d0743066f;
mem[837] = 144'hf5ceffddf089ef990f4ff8ed0dedf5a0f74e;
mem[838] = 144'h051c06ecfeedf794f86df4c20b83f1090b07;
mem[839] = 144'h03680d6603a40d510c00f18ef8c10d1f019f;
mem[840] = 144'h0df20063fa12fc2d02a0fe3d0a19065ff0e8;
mem[841] = 144'h0ed000fcfe54f39ffc9209f1036d06660701;
mem[842] = 144'hf44f00da05ddfbd2f045fdf6f780ff7805d7;
mem[843] = 144'hf317faf60047facbf2c6fa4407a9fccafef6;
mem[844] = 144'hf98af3d90c12024400cef8010a8100210a31;
mem[845] = 144'hf3150554036d06f3ffcb0c2d077304e80042;
mem[846] = 144'hf812ffe7f596056afffcfcd50afefb81f8af;
mem[847] = 144'hffd2f351f39e08390f25fe51035604af0ff0;
mem[848] = 144'h06c80d2efb9e0323fd2508e3f6ad005bf942;
mem[849] = 144'h0702fc92feeaef2909e100c209b2084c0a30;
mem[850] = 144'h05200511033301360d81ff9102b9003cfa22;
mem[851] = 144'hf216f66000c10d0df68d0895019104ea0565;
mem[852] = 144'hfa8bfb3bf575ff5406ccf2320794f25ef996;
mem[853] = 144'hf534f568f7d80338f3d0f500fcbcfaa1f3ad;
mem[854] = 144'hf4ddf6db09b10363f6a402d6081af04e026a;
mem[855] = 144'h0b33fe7d0ef0f31df029f677fc0b026d079d;
mem[856] = 144'hf526fdf9f6daff3c090c0e99f64ffbfd0cd6;
mem[857] = 144'hf0d30a1704ddfb9c008c0af806910e4bf95e;
mem[858] = 144'h0c81091cf73afda8040c025a0a09f5f5fe36;
mem[859] = 144'h01a0fc76ffc000740213f1c2fcb4fba7f7be;
mem[860] = 144'hf43efacd0b1606cdf9230e11f37ff148fd7a;
mem[861] = 144'hffe6f26e08eb0939fbddf52b0e6304670ef1;
mem[862] = 144'h022cfea1027bf7060db2fb2efa3ef2190e07;
mem[863] = 144'hf5640a160ed0f546060df331fd9c077600cb;
mem[864] = 144'h04f9f501ffddf2a4f06a0f370939f75af42a;
mem[865] = 144'h04fffe6602c3fe09f2230441044df0c30688;
mem[866] = 144'hfb9cf357f237f0c30c58044d0d730c8df520;
mem[867] = 144'h0be006c2fd02020ff386fbb90f95fd39f467;
mem[868] = 144'h0f4603ed03d301210473fd21f1b802e50827;
mem[869] = 144'h0d1cfa6008390ecefe9601dbf0a7fa220c3e;
mem[870] = 144'hff62f446f1b3f20407bc0ac10214f60d07e4;
mem[871] = 144'h0ebaf8fa031701e3071707dbf1f9fa3b0cad;
mem[872] = 144'hf206f3c50cc7f2dffdf8fb6c0e3cf5a30124;
mem[873] = 144'h0eb4089804110865fdf5faab048200c7f50f;
mem[874] = 144'h07aa092a05340dea0bdcffd8f5280603f8bf;
mem[875] = 144'hf0b7064bf991f3f2f2230157f5300c1bf184;
mem[876] = 144'h0ce40d55f877f2bffcf70e72012cfea600d9;
mem[877] = 144'hfa820fd1fb170a4b002d0a4d0f76f24a0b93;
mem[878] = 144'hf65f0addfedcfa8f05c7021a006af5650759;
mem[879] = 144'hff3d02e5fd88f43ef35a054e0ee50604f2a6;
mem[880] = 144'h0703f47f0f5a06720ce50b3305fbef87fa4b;
mem[881] = 144'hf4770867ff590123f2640e120d69f5bc036f;
mem[882] = 144'hf66ef096f70bf2910ba8089c05ac061304a1;
mem[883] = 144'hfb17f2d4f96afff10371088600ebfe4bf1a7;
mem[884] = 144'hfbf607280deaf3a20f33049ef14c00a20789;
mem[885] = 144'hf523f2befce60a170a03055903b3f8dcf2f5;
mem[886] = 144'h0721fee804ecff7cfc040220055202240d0a;
mem[887] = 144'hf4c1066608a4fc27f648f1d7fae5f8840d96;
mem[888] = 144'h0bb6f1e207b005b10693057cf89308200aaf;
mem[889] = 144'h08a109e2f061f1e1f7d9fc35fae2fd2303c4;
mem[890] = 144'h08ab0122f7de06130845f0c7ff52f009fcbe;
mem[891] = 144'h0f4df176081afb090abcf546007ef7d4f466;
mem[892] = 144'hfff7f7a3fc28fe33f3c0040b0f7cfdddf3b8;
mem[893] = 144'hf6baffc4fc91f0fdff380ec10270efda0247;
mem[894] = 144'h09cbf670f2cb07c1f3d20ec2f31608ad050f;
mem[895] = 144'h000a0edf08c8fecc028bf8d8f8ea073f0306;
mem[896] = 144'h0b7a0a440791f7de089b0c670011fb7af763;
mem[897] = 144'hf0ee0076f3d607e6f7fcf189f13a0aa3064b;
mem[898] = 144'h06c5f5eff444fe1ffa1605d0fc8efef7fdf1;
mem[899] = 144'hf52e086b07810f1af4ffeff50c630950f9ed;
mem[900] = 144'hf3ff0420f99d0d8f0bc303a807fc0300006a;
mem[901] = 144'hf469ff080c0708c2fe31f2b5f08afa14f21e;
mem[902] = 144'hf9160dacf8850413f471fbd3f329ffba05cf;
mem[903] = 144'hfc0502b407830cb4f91afcd7f4a4f12f082a;
mem[904] = 144'hf7ec045a0d65f78df9aff885fd5b0f800e5a;
mem[905] = 144'hfc0f0ec40c8cf07703a90d97f027f941fbda;
mem[906] = 144'hfe4bf100f8310a08fd630647f66506e7fbe8;
mem[907] = 144'h04770c19055e08c905880928066c0df10a0d;
mem[908] = 144'h095ef162ff4ff2120763efd60d80f5b90105;
mem[909] = 144'hfca207b9f3c3fadd06a7f28300e7065ef067;
mem[910] = 144'h098a0a7607b4f4b9f960f39dfae30ce3f404;
mem[911] = 144'hfba3ffaa0d63fbf2f0c602180d8f038bf897;
mem[912] = 144'h0aff0cdbff67f0eaf567f691fd600dd1f24e;
mem[913] = 144'h072402190d3bf9ca0e2ffbd8f073f0fff18b;
mem[914] = 144'hfbc4f035066cf247fdbc010effdf01e1f886;
mem[915] = 144'h07bcf42c0ed5f3e20d8ff13e060c0a2df954;
mem[916] = 144'hf1f5043df3fb070bf058fee60771ff56f115;
mem[917] = 144'h0270f14e051afc89efc0fe19f34bf02f02de;
mem[918] = 144'hfc870477fa84fe4ffa60f4570907fb54f179;
mem[919] = 144'h082f037205fafe2cf814f9b8f844f095f72d;
mem[920] = 144'h0977011e08980a8605adf978f5fff7f2f20d;
mem[921] = 144'hf5b0f3dd08c008e9fa15000c011c0353044d;
mem[922] = 144'h0a4e03b10f750e60ffe40b7af840fd67f853;
mem[923] = 144'h0f59f4890356f76f0fc00370007bfebff912;
mem[924] = 144'hf5f5fe87efd5f4a70c06fd580325f7610798;
mem[925] = 144'h089ff67903b5010d060a0da2f38306a103d3;
mem[926] = 144'h01f3fd65f844f80bf3f304e6fbdbf0bcfd11;
mem[927] = 144'hfb77f4cbfaf509f504d40d32f2f5ff67f12f;
mem[928] = 144'h069ff771072b0759ff54fe1100adfcadf726;
mem[929] = 144'hfcb3fc910a2a0c8b0398047d0c1804ecfef7;
mem[930] = 144'h063afbf7094f071fffc9f6fe00b907ee0b7b;
mem[931] = 144'h046b0970f5dc0dcd08490f790f36f53cfaaa;
mem[932] = 144'h0e0ff75003790164fcf5f24700f00906fe35;
mem[933] = 144'hf8870d28f5ee0831fbd90f450878f088fbd3;
mem[934] = 144'h05a8fbcbf001068309b3fefa0a86f48d08e0;
mem[935] = 144'h0ee7f959005b05a5093f0d8ff2c7fc79ffb3;
mem[936] = 144'h0b3903b9fd0902c0f55dfcc4faf9ffa2f329;
mem[937] = 144'hff56ef980e11f4e2f0d40de8f461f8edfa15;
mem[938] = 144'hf7240beef6aefa580428fa16047fffa5f291;
mem[939] = 144'h0eb8f1270731fc1ff0b00da70b99fd72f738;
mem[940] = 144'h06670bb7fb790713f0650d3af8620cd8084e;
mem[941] = 144'h0a2a0e4f0b780e9f0cb10bc2fd000c18f76a;
mem[942] = 144'h040504ee053b0baaf40efd640541fa6d01c2;
mem[943] = 144'hfeb9fecbf12c00f503cf01a7f5d7f400f411;
mem[944] = 144'hf614f8d5081206ed0732f0ac0aabf40e018a;
mem[945] = 144'hf1fefa92083af6ff0a7bf3b10bbff3310ae1;
mem[946] = 144'hf37d0147ef9b0a890cdd0d1109370a24eecb;
mem[947] = 144'h029df44df158ffea07660e1f0bed03ddffd4;
mem[948] = 144'h0383f6b40295ff6ff05af201068f066d09c6;
mem[949] = 144'h0e5d07a6f7eef5f2fcdb05cd0686fa550dfc;
mem[950] = 144'hf6ed0d23f190011b0848f564fc27efee0ae8;
mem[951] = 144'h089d0ea00b2efc9a08baf31cf57ffd5afc49;
mem[952] = 144'hfd81fc1209e10d93f439fdfef66ff7a70e70;
mem[953] = 144'h02ac074509d9fa68fd15fb8cf3e6ff6507b2;
mem[954] = 144'hf21efa5c0d390634f434f65bfce1f452f979;
mem[955] = 144'h0f7ef063096d0045f6cc0f92f60f06e00252;
mem[956] = 144'h0e1a04d10eac05b70675fc7a0accf046fe8d;
mem[957] = 144'hf92b0440fe29faebfe1bf9dd04d109720c21;
mem[958] = 144'h0b520391faa2fee20d53f231062df30f025e;
mem[959] = 144'hf9cf02df07d5f22cf19e03a90aa90ed1048f;
mem[960] = 144'h0c810e26012bf098fc14ffb8fbe0f7bb0392;
mem[961] = 144'hfea4efa6fffb0dadf0680124f51bf7770db8;
mem[962] = 144'h0d48fba5032a0119062afe1c0030f037f299;
mem[963] = 144'h0aedf24af2d0f5aaf4bdf459f7fffa1df9cf;
mem[964] = 144'hfffd01c70679fb4202990bcef4e0fdf7fc71;
mem[965] = 144'h048ef756fd770b780c2601730c3ff0e5ffeb;
mem[966] = 144'h0496028b0be90879f668fdb00014f18c0df3;
mem[967] = 144'h077c0d220bb3f5d4f21fffef06fbff95fa05;
mem[968] = 144'hefcbfe33f68c072e0a99f94afc9ffb0cff33;
mem[969] = 144'hfa62021c00d3088dff4af2ee08410f6a019f;
mem[970] = 144'h0279f707fd3fff260463f7b3fc9f033b0aaf;
mem[971] = 144'hf2edf853fe0e01ecf8eb0f5c03e9fec80c43;
mem[972] = 144'hfd750d7c01c3f3550db10878fc9bf0ee02b5;
mem[973] = 144'hfbfef9ee0523f7290eeb0f0b06d602a6fcf5;
mem[974] = 144'hf33605bcfe99f3f401c4081b02520a5bfd2e;
mem[975] = 144'h09de00cff42203c50ef1f5daf59a045d0572;
mem[976] = 144'h0d250cbef1230d93ff3e04d0f9b0ff890366;
mem[977] = 144'hfb760b540ef1fdb1f0a3fbf70855044effa7;
mem[978] = 144'hfe5e0017041bfcd6faadf315020ef9b5f465;
mem[979] = 144'hf6e2f59cf6ac0ec1061e09e604eafbd80af2;
mem[980] = 144'hf6bcf368f28cf3ebf562076f0b53ff1ffa23;
mem[981] = 144'h072ffce4027efd68f0ba0c58fbc600d701c0;
mem[982] = 144'hf5610064083ef8b600260ec2f3c6f45cfa81;
mem[983] = 144'h0c25f9f3f1c1ff8603fb072cfc38fb72fb66;
mem[984] = 144'h0e640d21f80cfe3503fbf2c8faa00260055d;
mem[985] = 144'h0b68f69bfd5cfc1bf2a70bbdfc76fc54ff04;
mem[986] = 144'hfc54080e06cdfb530744faf4fd31f742081b;
mem[987] = 144'h0bda06e5f0e1f5f60f1ef0bb0936fb9404ec;
mem[988] = 144'hfa0402e1ff47f0f5022ef09e0015024b0995;
mem[989] = 144'hefc701eff7a60e020afbf741f8a6f375fc48;
mem[990] = 144'hefecf80e0658f03cfa0dfd6f0b24ffac099d;
mem[991] = 144'h0d0c0fa00fba04a40e0808b30be502e3f3b5;
mem[992] = 144'hf130f78ef2fd001909b7f983f7db0d12f7e7;
mem[993] = 144'h063e0d87fa73fd0f0be408620a860689fde8;
mem[994] = 144'hf466f44e04960e200a9cfd07fa180cfe008a;
mem[995] = 144'h05ebfe81049efe0f0bd8091ff40f024af206;
mem[996] = 144'heff6fb1af209f5a1f3d90df900c00ceff257;
mem[997] = 144'hf7ff0962fbd2088efd57fdcf07db0c7df839;
mem[998] = 144'hfd3406660d970e53f8c404170b69f6e8f10e;
mem[999] = 144'h0639ef7906d4ff7bf29300450b6700f3f8fc;
mem[1000] = 144'hf1b2f8ddfa6509a6fb71f8990698f7d7fded;
mem[1001] = 144'h0c140c560cc1fd3d08f6f13bfb0a0a8304f9;
mem[1002] = 144'hfd99f02df8dd07d7f17b0a54f5d8f2a60d57;
mem[1003] = 144'hf4b1028402e4012bf318fd75f7c40119feff;
mem[1004] = 144'h09ed016f0a1f0c32f5ea061cf3aeefdff877;
mem[1005] = 144'hefa30c7b0c2900b0099b0c0ef83008eaf9c5;
mem[1006] = 144'hf052f309fe15f2690a35f680fbe6049500d1;
mem[1007] = 144'h0756f5ed0b400e9cf5c5f873f1d3f3200ce8;
mem[1008] = 144'hf32af0f505fff8980308fffcf30ef8a5fd98;
mem[1009] = 144'h04d40d97fd4c0e59ffb9f183080ef50ff2b5;
mem[1010] = 144'hf0840561035507fc0ab700f6f80df1c70a09;
mem[1011] = 144'h0e3c06e0f1b508b6f12e049af685fbf20d16;
mem[1012] = 144'h0b69f7c3085efffa07a6fd6b024ff0be0588;
mem[1013] = 144'hfb1a03bcf6f4f39e0729fdb3f97002adf4dd;
mem[1014] = 144'hf6fefaa203d3f210027b02bf0af3f363f285;
mem[1015] = 144'hfba8f6130a5ff1270a66f7360e2808350d90;
mem[1016] = 144'hfa3604d1f607f1500262fb6903cf07fc0d84;
mem[1017] = 144'h037d0807f0b3f550018efc75f4f9fb4a042d;
mem[1018] = 144'h051d0a49f12f0ce2f653fc7f0cb10655fb26;
mem[1019] = 144'hfe000119f588ff48f61708be0317faac0753;
mem[1020] = 144'hfa2c0e9c0b5df9fc06bf0c2103c709c20add;
mem[1021] = 144'h0e0defa80269f59f04ddf6ecf83f082a08de;
mem[1022] = 144'h0ea90547071c0f59fa4d0d4df552ff4c0cf4;
mem[1023] = 144'hfdb6fba8f04e030309fc012b00d60fb80e40;
mem[1024] = 144'h0c410e38f1b50217fe0a042bf1dbf15df066;
mem[1025] = 144'h0c28f138074d0684006def380f460c16efe7;
mem[1026] = 144'h0b800efcf68d04abf1d90d8a03b20c13fd88;
mem[1027] = 144'hf49f0a5f0785fb0403a80e8304cb0efb0cdc;
mem[1028] = 144'h0d8efa40088703a70b3e0a6a093a06f0f061;
mem[1029] = 144'hf7f1f3ec0bffeffcf6530572f96d015a06de;
mem[1030] = 144'h0da3fa320696097ef8b207a9fc0906c6f8b5;
mem[1031] = 144'h0526f57002b6f858f7d404a400d806fc0980;
mem[1032] = 144'h09acfca2feb90227f78df61f0687f3300642;
mem[1033] = 144'hf9ad03aaf0d70d270263f1dafa5a07dd0d94;
mem[1034] = 144'h09f60dd20dc4f54ffb8c03770756f13cfa89;
mem[1035] = 144'hf6fcf551feb8ff41f059f5cefd42fc9af9a2;
mem[1036] = 144'hf9f00506fb0306a2f39707810d660d05effa;
mem[1037] = 144'h081b0b85f496002ef28af58408a7f458f7c0;
mem[1038] = 144'h0bcfef59fc1afa320aee02ef0b08064907fe;
mem[1039] = 144'hf4d5045b070ef8b0f627f5570ab6f4a2fd26;
mem[1040] = 144'hf38a0fb3f5f20b14fcc7f26dfdc507faf069;
mem[1041] = 144'hf929f166f0dc05cf06b50884f1180327fbce;
mem[1042] = 144'h004cf406f54af7c30bfeff1ef5a8f158fb3b;
mem[1043] = 144'h0999f1fbf27c0ad1fbddf0a3f4ed0b34f31e;
mem[1044] = 144'h00d9049c0d8cf3edfd260fcf0536f343fa4a;
mem[1045] = 144'h0515fd2402aa04900ab3008df8dd093af5d5;
mem[1046] = 144'h099f0ad0fed5f60f0f850a31f4ff06a406fe;
mem[1047] = 144'hf5e10845f15df84803f7f5f5f3dcf3c1fd8f;
mem[1048] = 144'h0b20fd5f059df74a06e000d4fb97f4f70516;
mem[1049] = 144'hf74def5dfaf009730f310dcdf3fdf1d7fa6e;
mem[1050] = 144'h078d08b105c9036e0be8fa8801a8fc560102;
mem[1051] = 144'hfb4f0e94067f02560dfc025cf0a3fcb20de6;
mem[1052] = 144'hfd900c9efb0a0bc0fa81f626f8d808a5ef0a;
mem[1053] = 144'h0bd60300fedcf890f14204d5056c0ab30052;
mem[1054] = 144'h0998087cfe1cfc2ff3a4f3ec032cf7a30e90;
mem[1055] = 144'hfffdf42e017bf89c023ff70ff70a02a6f2b2;
mem[1056] = 144'h0d7dfb8b0703fc2d0139f3f2fe8fef79077a;
mem[1057] = 144'h030e0690f16104e1eff50d47fb38f126fc36;
mem[1058] = 144'hfcd2fbc606cc08e7fea7f15cfabcf6c0f3a5;
mem[1059] = 144'h04aa077605cb0ba2f1a005440c61085ef641;
mem[1060] = 144'hf68ef68eff800a82f4cb00fc0909002cf91b;
mem[1061] = 144'hf5c40902f5130296f386f487fb32f4e703d3;
mem[1062] = 144'h0219f60efcd8ff34f6440745faf3009bf018;
mem[1063] = 144'h0f57040ff2000d3ff9f303d4057e02b60219;
mem[1064] = 144'h0c1efc8afc320036f2c805e8efedf40b04c1;
mem[1065] = 144'h09f3fd29ffdcf8810a11fbf30b3101eb083f;
mem[1066] = 144'hf64f0ccb0800fa10fcbdf694fb330ceff4f3;
mem[1067] = 144'hff70f7b6023ef7fdf54afae409eb0047f45d;
mem[1068] = 144'h0b86fe30faadef47f7d7f923047dfdea09a8;
mem[1069] = 144'hf9800b1e0a4cef5201ba04b7fb18f657013a;
mem[1070] = 144'hfcf9097b024005f60d97f7dbf8b70950fe9c;
mem[1071] = 144'h066e0e8af9e3feeff7d60a2b0dea03590a97;
mem[1072] = 144'hf515f649ff6fff3ffea30da50a4103940c74;
mem[1073] = 144'h0fb5023ef5410119f047fda0fa6300c209dd;
mem[1074] = 144'hfc0801eb0670f04c0deef1daf4b6faad049d;
mem[1075] = 144'hf5c5f044fedbfaa5f041f33ef4c1ff55ff78;
mem[1076] = 144'h055ff7b4ff3f0a62fe8af6350a15f37402b3;
mem[1077] = 144'hf16809e7ffe60f260ad90a9a0a1f06150422;
mem[1078] = 144'h0b6805a9f9e2f019090c00c50985fdd0f1a5;
mem[1079] = 144'h04fd0c8608d1fd790e32f4e201d7fd41fb6f;
mem[1080] = 144'h0c7b0f0ffffaf9bcfd45043c02f2056e00e0;
mem[1081] = 144'h045808affa5b09600daa042007c1f2210d1a;
mem[1082] = 144'hf70d05430c75fa89f1b20479fc6907f0fc09;
mem[1083] = 144'h017f0be1f4aaf34ef485f38af01a0f89075d;
mem[1084] = 144'hfd07febb07e00ba8030bfcdeff95f270fd9d;
mem[1085] = 144'h0870f7adf1d703980ca70b07fcdb0a15fae2;
mem[1086] = 144'h04bbfeb90301f514f64a058efcdaf85d0bd5;
mem[1087] = 144'h042c08fe09aff775ffa4f8a3f31d01f60796;
mem[1088] = 144'hf9d3035b0bd90f19026df3e8f934ff930a31;
mem[1089] = 144'hf4b2f869fd2dff1c0443009d044cf88cfe2e;
mem[1090] = 144'hff77058c11f2f56c0996ff93fe90f255f6fe;
mem[1091] = 144'h0d3d0e26f3420f830f63f0700b68f05dfac3;
mem[1092] = 144'h0603f766f39905b4f4b20fdb0bf80841078a;
mem[1093] = 144'hfed5f51a0afffee1f4b802bd039905970c43;
mem[1094] = 144'h05e5f9c7fd7efcfc00f2fd440127f9a60d12;
mem[1095] = 144'h037c04f401a20452f157f9aeffd00050f749;
mem[1096] = 144'h073ef74c07faf7830b22fc300058ff6bf1d5;
mem[1097] = 144'h0006ff1408220094f3e00650021e0afdf923;
mem[1098] = 144'h0144fca205dbf879f042fbac029df0eaf623;
mem[1099] = 144'h06df0699fff2f08e04e4f7b101dc00ab0375;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule