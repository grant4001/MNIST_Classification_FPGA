`timescale 1ns/1ns

module wt_mem6 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'hef36f76603d5fa10feaff4ce07dbf26bfc3f;
mem[1] = 144'heebd04b5f1f9f8ddf84ff4aef35d076cf00d;
mem[2] = 144'h08adfa64f79c069d07600a4c025eff6809a0;
mem[3] = 144'hf1a705e108f0023103d4f79fff2c0bba0533;
mem[4] = 144'hee82fbc8f80e0415ff1e0a4df4d50b32f5c0;
mem[5] = 144'h0467f596012f0c34eee9f7c3fe5000fef004;
mem[6] = 144'hf681fcb205fef216fd0df8cc018b037d0329;
mem[7] = 144'hf7adfc150762f51f0ac7fb690889fac6087e;
mem[8] = 144'h0544002b0a0eff91edd3fd980b58f0ce092f;
mem[9] = 144'hf87af45e0a95fc390410f230f00af8f80db6;
mem[10] = 144'h008104b704a0fe350719ffa404b6f723fa24;
mem[11] = 144'h04bd03f5f43f06a4f1a2f5d0fc060be2075a;
mem[12] = 144'hfeb5f920fbae0849f69af8c7ff7ffad9fe5d;
mem[13] = 144'hf88509900c5a07adfdd4fbad066401f8ef6b;
mem[14] = 144'hf2c001cffc09edff0b450de4f0bcf8dc0c2e;
mem[15] = 144'hfe79f1dafd7a0ae9fa7efb460251ef990db8;
mem[16] = 144'heb81fe91f3f909adfd00fe00f0a400c5064a;
mem[17] = 144'hfaaef967ea1f05620129f8c50988fe780051;
mem[18] = 144'hf088f3c7fbc1051ef532fb7df462f644f6ea;
mem[19] = 144'hf5fcf70c00fc0255fe95ffc202880901ef6c;
mem[20] = 144'hf515f844f1b5f861f80ef3f9067ff7ffeedc;
mem[21] = 144'hf7cafe3df301fc8af448ed62edb7f412097b;
mem[22] = 144'hefb7ffea07c0fa73ec5ef3c5efffff59fb0b;
mem[23] = 144'h06d8f7e2fd08024bf050f05ff40902abf155;
mem[24] = 144'heed7fd3ef99ef6d90908fd30ffadfee20383;
mem[25] = 144'hfb66fc9afb65f383048f0034f4adf8bc09ff;
mem[26] = 144'hfb1af2c0f544eeecf286f89d059400ecfabb;
mem[27] = 144'h07c40ac9f4dbfa58f6ebf9fe05e9f2aef79f;
mem[28] = 144'h0da9ff690b0af1aef190fca8ff190bc4074f;
mem[29] = 144'h06adf1f0f03f01ac0dc0fd8f07bd09d7f94c;
mem[30] = 144'hf7d30b80041906f8ed1306d6f90fefab0250;
mem[31] = 144'hed54fe8ffe33ea24ed8de991fde001bce968;
mem[32] = 144'hf772f99bf085042cf687ff6ff142f73bf557;
mem[33] = 144'hf2c70a61fa2cf76cf56703fbf74ef754f24b;
mem[34] = 144'hfcf4f81205a3f54ffcd1055801d106990799;
mem[35] = 144'h0a9005e40262ed48eedfeab0ebaee8c10425;
mem[36] = 144'hf798f93700cbf69103b8fa6cf326f483fb49;
mem[37] = 144'h08d708affb7af263f3b908a2096aefd8fcae;
mem[38] = 144'hfb2f03c1020ff1e4f6dcfdf2eee801d802fb;
mem[39] = 144'hff2502b3f9b1f1690093011eed7af31afe20;
mem[40] = 144'h0283fa4c01ca0b8f063ff19302d6082d0bc2;
mem[41] = 144'h05c5f25eef3102c60e11f06bf096fe30f32f;
mem[42] = 144'hf6e6faa8f3bfedbbf5ee07fef8f7f77b06ff;
mem[43] = 144'hf8ca0b64098feeb2ef4bf8c60497f10a077b;
mem[44] = 144'hef81f5fafa2df65003e501a5f440fa98ecc9;
mem[45] = 144'h0186e999f742f7c105b0f3fa0335eaf4ecad;
mem[46] = 144'hf9af0cfefa8ef9f3f74b055bf729f3f4042e;
mem[47] = 144'hf69502d4f837fddff30206b602f8f321fc69;
mem[48] = 144'h05ecf3a6f3080052f37fed58fd1afc98f203;
mem[49] = 144'h0a21ee61eeb9fb9cff8c0009f718f2e5f72c;
mem[50] = 144'hfcdff370f523014afaa3f82af9750b88f7f7;
mem[51] = 144'hfff1fe50fd39fec2fe07fd47f303f28cf3f4;
mem[52] = 144'hfbf60a8e07e2fa59fedbfc85fec6feaff7d1;
mem[53] = 144'h03c9f27108f005b4fc7eeda30028f17ff7e8;
mem[54] = 144'hf245089702b5f0bef501ef10f904062506ad;
mem[55] = 144'h0b37f647f177022f0637fd0af0950750f4cf;
mem[56] = 144'h0ddf0320f77202e7fac00599f3430dd0ff62;
mem[57] = 144'hff0eff24f75ff1d4080604040c37f19cf35b;
mem[58] = 144'hf02f004af3e2f166facff40d0ccbfb06fa83;
mem[59] = 144'hf96def45f7420c2f039cf1850a78090bf80c;
mem[60] = 144'hfc650609f76501e8f96cef4cf07c07edf200;
mem[61] = 144'h04bef1f6f07af6e70b47fad802b703560064;
mem[62] = 144'hfdcf003c00c405f3008f095cedd307a00aab;
mem[63] = 144'hf02105fd01b0fb5b0ae802adf260ee00f5fc;
mem[64] = 144'h09a609b0f485f9ea0a1a066ced19f81dfcf1;
mem[65] = 144'hfbb300aefeeff188ff4c039af338f617f564;
mem[66] = 144'h06e4f222002d0564f2db0229f2af03310c45;
mem[67] = 144'h070afd94f9c1fecc0aba05440d720b280f4e;
mem[68] = 144'hf9d7f0480166098b07b5f95807dd0641fedc;
mem[69] = 144'h0db3f3e1f89a0e47073bfa840fb403ee0348;
mem[70] = 144'hf7c9f86ef70ef9b7fe92f044fcbe06da08c3;
mem[71] = 144'h0968f59c033ffbe7f9d9f4f1f1250aaa0875;
mem[72] = 144'hffb2f60d0ce0f61008c902faf911f75c0fbf;
mem[73] = 144'hfec3f9850413f2bd0be5f8e505eff7ce085c;
mem[74] = 144'h05e9feeffbb60bfafd200e9e0eb3f717feef;
mem[75] = 144'h02b20115f997f6e501b50369ff5df05605ee;
mem[76] = 144'hf0f0f1aef4b10bbefc9a0d32f87a0f4ef318;
mem[77] = 144'h0c29f3150c560afbf5b9006009e1fda60716;
mem[78] = 144'h08f907a100fa0261f147fc70f6cef4220502;
mem[79] = 144'hf9a50b750ea00d1703ef0ce2fde40ea30a2a;
mem[80] = 144'hfcf4f32505a501c0ff89f7fff0b2f4cff341;
mem[81] = 144'h0e4a048100daf826f4310ad0f7c30cfdf79d;
mem[82] = 144'h0fd9fae0ff8bf1ea0f56fe0df69ff0c3054f;
mem[83] = 144'h090a052af94e040704eefde4fbf007bbf96f;
mem[84] = 144'hfaa00818f5410046f88ffdf30ba502c50c21;
mem[85] = 144'hfd5ffc51f7fb014600b3f652fc48f928f1cf;
mem[86] = 144'hf3970992f93bf7ee09a3fb9df5bf0cb2fe36;
mem[87] = 144'hf692f11dfbd70e02fbc70ec301d4f1d8fbbc;
mem[88] = 144'h0aa10033f362f7abfe80fa15ff2afe910366;
mem[89] = 144'hf73e075df7880faef10efe54fba4f13f050f;
mem[90] = 144'hf55a06570acafea9f174f946f25200da000b;
mem[91] = 144'h0b13f005f58104380017044a043a04160d3d;
mem[92] = 144'h091f07f7f2e6007df82af0f30fa0fc34f2e1;
mem[93] = 144'h0560fdcc0da700080854f2230e5bf2d60af3;
mem[94] = 144'hfbccf0d4f9df035cf30af70703a4f78e0b5f;
mem[95] = 144'h03a80b0cf06c0fabfe09fadef77ff3c8081c;
mem[96] = 144'hf92d0bc00e4cfc07fd2ff7420d69f2d8058f;
mem[97] = 144'hf8550720fae30c0ff89f08400a680d35f99e;
mem[98] = 144'hf299f59c0b59fc1f04aff0dc01e0fc67f3d9;
mem[99] = 144'h0e05fa4dfd8cffff0bcff0f00fa705270e2a;
mem[100] = 144'h0dad065a0cc8f3c5f7d005c2f0b40c3f0737;
mem[101] = 144'h09da0eba0df7017c048ef24afad8f42cfd5e;
mem[102] = 144'h032af9f709a9f14ef39205dd0baaf3a7f383;
mem[103] = 144'h04790c03010c0039fe72fed70f22fc3ef587;
mem[104] = 144'h0779f7160261087900a50c2afe450e120dad;
mem[105] = 144'h0e5607b70556f28007c10c2d0499fbabf1f8;
mem[106] = 144'hf916fbeb0f9f04b10b180c3ff60f05cefc2f;
mem[107] = 144'hf7a5fd8ff0c507e00b2afc860929f641fa99;
mem[108] = 144'h03fe0dba001f0f050adf08f30df50f70f64c;
mem[109] = 144'h0d0c0d0dfec1094e0955f24a0922034d066e;
mem[110] = 144'hf8e5feb3fd02fadaf50703effab20458022b;
mem[111] = 144'h0dc509e0fda00abbfadef487093bfffffc61;
mem[112] = 144'hf47bfd9403310682f6edfdcbf6280032fa79;
mem[113] = 144'h0466fc4f02d1f26df0bdfe5df8140186f300;
mem[114] = 144'hfefbf7df0ee9ff7ff910f19704f8f19c06d6;
mem[115] = 144'hf185031c016909560b84fe280163f36df55e;
mem[116] = 144'hfef9fb6702170c07f549f8170b2f0e8702a3;
mem[117] = 144'hfe0cf745f4cff95407a60d2a0671081bff00;
mem[118] = 144'h0ef306d30c54f658fc45fcb90c52fddf0fba;
mem[119] = 144'h062f0f3afa01fbf10d5af29b069b00acffc2;
mem[120] = 144'h002effc2f7b2effd0e660efa0e760a300bf1;
mem[121] = 144'h035c0ed8f8ea0995062d097502af050ef3ae;
mem[122] = 144'h021c05e0f65f0fc809bff479eff507c00cf8;
mem[123] = 144'hfcebf1dcf80af4b3f6f9f5f104a909860c38;
mem[124] = 144'h01e6f19efe0a04e70ffaf596007af28101b0;
mem[125] = 144'h02470b8a036ef4f8f36ffdd80c47f9b5f219;
mem[126] = 144'hf156f438fe85f6000c800cae0fb9f0040a17;
mem[127] = 144'h0b8df21ff703f3b9f8e1078c0b50f52efa8b;
mem[128] = 144'h0e62f48a087efb620b43047205070c250b5f;
mem[129] = 144'hf21cf7a404b0f774f3d2f675f3c00b11012b;
mem[130] = 144'hf3000719085208c70bc6f77a0e0f0610fe26;
mem[131] = 144'h0986f69cf3eb0683085bfeba02050a8af009;
mem[132] = 144'heff305400b0cf689036d0be809d80b73f338;
mem[133] = 144'h0868f922f749083f0bcf0e6d03ae049df911;
mem[134] = 144'h07de0d2c09fcf95e0acdf79400490ae7059b;
mem[135] = 144'hf3200299f62302ca05dc0b700ef50a970485;
mem[136] = 144'h0f06fdc9072cf1aaf5430d4902e3fd25f2d2;
mem[137] = 144'h0a5cf1ec0d9df5030bdcf021f03b076d094f;
mem[138] = 144'hfcd1fd4e071bf2be007608f20bf90a2f04b7;
mem[139] = 144'h06ab0402044df171fa25f56df62ef9ff0be4;
mem[140] = 144'h0c93f45c0afcfb9dfd2605ed0c2efcea095a;
mem[141] = 144'h0ecf0893fa690503085ff3fbfb22ff1df81a;
mem[142] = 144'h043907f90cdb0d83ffaffd15ff88f00afa0e;
mem[143] = 144'hf0d00689f9e8ff27f1d3f267f2a5fea80269;
mem[144] = 144'hfd7cfd4604fe074e08640c03f4c0f11c01b1;
mem[145] = 144'hfeb60d230ea80004f8dff05106d7f8e0ffa4;
mem[146] = 144'h071df937f7bdf4b9f0f6f3e4f14900a20457;
mem[147] = 144'hfee3f611f42c0238f549f055f5effe8e0c1c;
mem[148] = 144'h0738f2e90f38f95703ae0128015efa40f0b3;
mem[149] = 144'hf03e07050211f3b30bb1fb750b32007bf8a3;
mem[150] = 144'hf3720673050f0f89fdb00e9df74d0426fe25;
mem[151] = 144'h0772fb9d0b7ff277092af0b20cb90d7cfad1;
mem[152] = 144'hf1a1effd03f30a1b05f9fb40ffb106ccf900;
mem[153] = 144'hf4bf0a8c06b40eb7f7a1f10df334f263fd7f;
mem[154] = 144'hf37ef00e0f8cfd1cf6d7f1f50b770d490b0e;
mem[155] = 144'h09700632f315f5fc056209fdfe8c030ef30e;
mem[156] = 144'h00e3f5a7f1250c7dff0df5c3f6caf56e0088;
mem[157] = 144'hfbf6f1710406f237fe8b057b0cc3fab8f116;
mem[158] = 144'h07720841f891f999f9d2039b0af40fea016b;
mem[159] = 144'hf892fa8609c20b980964023efec60f1bfa00;
mem[160] = 144'h0ca8fdc8f91bf87b084ef4bbf72102db0b37;
mem[161] = 144'hf402fdef08fd0e77086d02280a69f7ce07e3;
mem[162] = 144'h0cfbf77b056eff6c084803f7f52cf23f048f;
mem[163] = 144'hf8bff6a4f73bf4e8f26e02eef6b304c90b2c;
mem[164] = 144'hfca50a53097bf94e0dae0d32fdd0053cf2b2;
mem[165] = 144'h0fbcf469052cf522f71ef2d80e1e0612026d;
mem[166] = 144'hf562f2910f930ef30f7cf7e20d7d0a0bf4c7;
mem[167] = 144'h0f040d00fe57fd5f05180c44025d01040fb8;
mem[168] = 144'hf33af60afe73f426fb4bf3d7f6f3f0c8f189;
mem[169] = 144'h02d50348ff0909860a3e01360acef51efba6;
mem[170] = 144'h0afb0e090ef302630e38efccf0760b3a0466;
mem[171] = 144'hf83b0ab0077bf187fd5608acf9aef0fdff42;
mem[172] = 144'h05b80b63f27906d30c46f7690d46ff36fad5;
mem[173] = 144'h00700d0d027a04b4f362f26d05b804f0f273;
mem[174] = 144'hf179f7c2fa210e1005840f80096507760e56;
mem[175] = 144'h071cff0efef40028fffb0351f8750f1905e4;
mem[176] = 144'h08b7f635040af734f7b40edbf667fd440c8c;
mem[177] = 144'hf16c05f909a30070f25d01ae0ed108e30a1a;
mem[178] = 144'hf2b2f45b082af24c0c70ff36fde0fcf305a6;
mem[179] = 144'hf15b06a9f36704040025f9a5ff7e0cdcfa9d;
mem[180] = 144'hf0affd7f01bb0c030ea9fee7033b0ceefe90;
mem[181] = 144'hf23b0adff8d20f4bf9680c610f4cfe0c0108;
mem[182] = 144'hfa44000b0572fffefb9ff124f65af244f9e5;
mem[183] = 144'h0827043001a507d1f19a09b406c5feed0bfe;
mem[184] = 144'h07ab081208c9f9f9f275f78304a10a98f494;
mem[185] = 144'h0806fbe1fd13f3c0095200c6f4b80b46086a;
mem[186] = 144'hff330a78f298089ff454f9b0f01c0099f4b0;
mem[187] = 144'h03ecfc93f7aef53d010e032ef0cc02c0f020;
mem[188] = 144'h0e73fb8a0f5a00e30a7df59e0cb8f263f83e;
mem[189] = 144'hf5fbf9d4f04c002df44c061c0b2ef109096a;
mem[190] = 144'hf2c20e940483f78a05f805b2f88c0b370e6d;
mem[191] = 144'hf355f6b106c506bb0cf1f4cd0d16fc3c0430;
mem[192] = 144'h0d73f20805ba0f7302ebfadb08ce0ce6f56b;
mem[193] = 144'h0c33f1e0f27406de042408a502ec0320f1be;
mem[194] = 144'h009af6fd02ba091103b5f375fa62fdb3f1c4;
mem[195] = 144'h092bf80cf2f00d93f2f50a66f6fff382f31e;
mem[196] = 144'h0465f3400bf0f52609a8fbf0fab605eef606;
mem[197] = 144'hf565085c0098f202fcf4fc170cd6f57ffb4f;
mem[198] = 144'hf2b008b1f66302c00887f863056a0f3c00ff;
mem[199] = 144'hf68cfee605dd019ff1e7fc4e0aef00380e17;
mem[200] = 144'hf2ecfa14faa9f66af955ff61fada0d9907d9;
mem[201] = 144'hf3e90a60084e0bd9098af76df39c0cab097a;
mem[202] = 144'hfc3e0bb4f234f9f70477f769fa65f582f38e;
mem[203] = 144'h032cf130050e01e8052ef9c6fa140f51fef8;
mem[204] = 144'h0750019ff0fef1ed018c0103f3c8f0a80142;
mem[205] = 144'h0767f5d3f066fa6afc97f77405200bd9f1bb;
mem[206] = 144'h03daf7e5093ef831f0a2f3990acdf999f171;
mem[207] = 144'hf9b9f4aa08590e66073d027e0b6c065702f8;
mem[208] = 144'h01e80f23f5f6080aff2003adfb60fc1bfd92;
mem[209] = 144'h02860b7efda5048dfbf7047c0456f7960e9e;
mem[210] = 144'h01740a140a11fc8c06f8fdb1f2d504fff6ec;
mem[211] = 144'h0c8af896f5fa0f5bfde80d470dbf03320409;
mem[212] = 144'hfdd4f31af88e0721039a062b08bb0ff2f263;
mem[213] = 144'h005609adf6c70805f5fbf4e4f0fc0e5b014e;
mem[214] = 144'h0841ffeef4970742052a09cdfee406e6fdbf;
mem[215] = 144'hf55b0c270906f486f65404c805cc0dd60e34;
mem[216] = 144'h0402fafaf4b3f58a07e30d2605c2f0f4fc90;
mem[217] = 144'h0f62f8d9f9950ba9f2cbfbc200670c52fcb8;
mem[218] = 144'hf6bc0b55feeefa3bfcc7fe9f0983013ef9cd;
mem[219] = 144'h0bcefff9f9e3055f002d03740e22f148ff35;
mem[220] = 144'hfa8a0a35f7130efa0740faf404b101baf2dc;
mem[221] = 144'hfd5204b20226fe13f02803d4045f0299041d;
mem[222] = 144'hfef70c230c31f7f60fbafe50fe3cf4ea0721;
mem[223] = 144'h07ecfd66f40dfc6806140fa0f4c8f933f666;
mem[224] = 144'h08b00790fac1091001f5ff7404d9f01608e9;
mem[225] = 144'hf7310c6bfc500055fa80071f0ed1fd2cf1a8;
mem[226] = 144'h05ecfc1a0da8f78efed70cdc09eef6fdf560;
mem[227] = 144'h08d2ff6a05df0724f9fbf88ef8e2f086fcd0;
mem[228] = 144'h02eff3670e1d09c70c6d0838f318fffbfa87;
mem[229] = 144'h08ee0cc90219fdd8f639048af2c7f0aff2e8;
mem[230] = 144'h007df1dff6700fdbf47c097d0af50eed0c86;
mem[231] = 144'h0d25f5bd0995f6390092faf1f532f22af0bd;
mem[232] = 144'hff64058103f7f5dc091df8e20ccdfe3a0662;
mem[233] = 144'hf231f2f80e3cfe9804410525fd53f8abfc4c;
mem[234] = 144'h026900ae0572f5e0f0ccf8a401020c9efab9;
mem[235] = 144'h076bff32f7fbf74e0750fe75f7b1f344f06d;
mem[236] = 144'hf9ef030a0d61f03209a6f566000afd630276;
mem[237] = 144'h002f09b9f63bfd45f21d034efd6b0ac6080c;
mem[238] = 144'hfe08ff23f127f558f65e09f0fcee0188f855;
mem[239] = 144'h0e68086b037ff585f46bf3b10d2cf633ff36;
mem[240] = 144'hf1c8018d0f39f676fd47fbe9f17ffec8f9e8;
mem[241] = 144'h06f30edd07d1f367028001da0221f4f10946;
mem[242] = 144'hf995054b0431f2650839021bfcc9f2950dac;
mem[243] = 144'h0ac5f70b0152f600fc22f9780e7ff2eb0dae;
mem[244] = 144'h03c503cc0fb007bd009a0d12fe76f8bbf745;
mem[245] = 144'hfb7b0c37fb78f44ff48ef118fb87023df8f9;
mem[246] = 144'hf54c0531f32a0e71f317f40ff0cffb04f4b9;
mem[247] = 144'hf89709660daa0e09f2c2f6f6f47ef4fffe93;
mem[248] = 144'hff7a0301f8a30e6c06aa0448fa4009c8f29e;
mem[249] = 144'hf6520295ff7ef12e0c3df3fb06040382f77a;
mem[250] = 144'hff0804c2f37bf4490153f20b0eaf01860735;
mem[251] = 144'hfde0038cf7000ebd0b22034d0257045af3a1;
mem[252] = 144'hf669f17609590f90fa37037f0ccff74cf4e8;
mem[253] = 144'hff4e0685fd7cf2d00fc8fc25043405ce0736;
mem[254] = 144'h0bfffb75066cf1d7f6a8f1b4fcdafdb60e1e;
mem[255] = 144'hf8020d6cf711ff75f962f18cf1a7f830f78b;
mem[256] = 144'h07c20cf2f4130750fa48052bf16906350fdb;
mem[257] = 144'h0de508ee0dd8fae50f16f699f212f54af942;
mem[258] = 144'h03210dcbf069f25cf012072b04ebfed1004c;
mem[259] = 144'hfadafb4b00950b6a0fc0f2ef09f60cf30c15;
mem[260] = 144'hfe5ff66e0d5b0958fed3f1fe08550630fac9;
mem[261] = 144'hf949f049ff81f1660b22f1eef36e0fb2ff88;
mem[262] = 144'h025ffcf203d3efeb0efaf418fe4902fd000a;
mem[263] = 144'hf5d70cf60634088702980af4fae6088c067a;
mem[264] = 144'hfd58fcfaf05001b3f2f102c0f981f2230506;
mem[265] = 144'hf71807ca0588f495f933ff7c06a209eafa72;
mem[266] = 144'hfff7f3acf0b7f56af90c0a62f351f9ef07dc;
mem[267] = 144'h0b2c0c7500ecf4f60cbf04060d28f9e60f1b;
mem[268] = 144'h02440805f2f3fc3f0c4401680956f1cff5a6;
mem[269] = 144'h082d0b670a58fa72f98a0df0f30af666f208;
mem[270] = 144'hfa7cf22306d50b13f4bd03cb0c17f4a403e3;
mem[271] = 144'hf852f9330103024c040df085053104fafe79;
mem[272] = 144'hf929f58d098703e8f999f97cf121f115f381;
mem[273] = 144'hfd5cf5d6ffe707230ae40d43f1800571ff15;
mem[274] = 144'hf61efd69f5a80d71f62a0f2701f00716054e;
mem[275] = 144'hf5e2042e0dfef3e50bc206fefaf3014a03cb;
mem[276] = 144'hf156fd4ef12e0654f7e0091103ca0fb701ad;
mem[277] = 144'hf4a30184fdc50ed30d4b00f5fc91f51f018c;
mem[278] = 144'hf69aefcc05bc0c41f483f216fd2cff3a071c;
mem[279] = 144'hfdb108fb06e108ad048cf28509c406bd0bfa;
mem[280] = 144'h0268094d0ef40879fd33fdaff2c7fa6cfc24;
mem[281] = 144'hf9f5f7bbfa0d0f76f80bf2990e9707c80044;
mem[282] = 144'h0001067df595f78e0dd50c580a0901e4fe41;
mem[283] = 144'hfd0306baff6a0372efc007b5f656f6040343;
mem[284] = 144'h099d06e9f9660a6b0ba9f76df4bdf01af4b6;
mem[285] = 144'h019af5860a96f2f3fc67efe1f4a2f14c0d42;
mem[286] = 144'h0266fb4ff34afa000cf90d0ffea9f9f6fce6;
mem[287] = 144'h08eff9df007ef9160cfcf9ef015608560cd5;
mem[288] = 144'hf08ffc8f09c20e6402b50202028ff22a018a;
mem[289] = 144'hfd8bf5760c0b04380edb0f6e0aff0c81fb2f;
mem[290] = 144'h04eb035df0d0f68af2ed02b3f00903950535;
mem[291] = 144'hfbff07fc045607ad0e4106eaf094049d0c9b;
mem[292] = 144'h06f609e302c008e80841f55feffdf6bb0efc;
mem[293] = 144'h0ce708c80dd2f74e08d10d31078d0010fd5c;
mem[294] = 144'hf4e10575fa3cf7a9fb380a8ef16d0a7f0746;
mem[295] = 144'h0d1409daf637018dfb5e0cbef00f06bcf404;
mem[296] = 144'h07e505eaf3a80b0e0d1b0a7ef66cf685fdd1;
mem[297] = 144'h003cfc6efc3dffbd01c6effafcecf6d70de6;
mem[298] = 144'hfa4f08f00ad9f808083bf2a305f1ffa5079f;
mem[299] = 144'h09eb0ee0f95df192febdf149f470f900f233;
mem[300] = 144'h04050390077b09c100100ac6f23d08ddeff7;
mem[301] = 144'hfc5af17bff1ff1f3f9790720fcfcfd0ff166;
mem[302] = 144'hfd0c02f8f772f452f5ddf1460a1708f2f9d6;
mem[303] = 144'h095a068cfa7a0ec8fd400365ff030adb0221;
mem[304] = 144'hf092f6e00bfb015dfdff055a053df906fefd;
mem[305] = 144'h03c4f94cfb230b44f657f9840c39023ff927;
mem[306] = 144'h06500f060de50e9ef52a000b04b10cb4f28b;
mem[307] = 144'hf82cffc006fef188f82103defad6f78cf6a8;
mem[308] = 144'h07acfa86fd78fba603090aa6f07afd43f743;
mem[309] = 144'hf8b3f2780e14fc3ff535f5500be3fcfd003b;
mem[310] = 144'h0314fe94f5a4f2c2f55802ba0d8cf22909d0;
mem[311] = 144'hf5ee03720c62062005390524f78505d7fa90;
mem[312] = 144'hf34d0eccf74aff57fd94f3900ef40c190956;
mem[313] = 144'hfc4f022500de0dcb0a61f6e700e7ff5bfb0c;
mem[314] = 144'hf394ffa7f59b068ff0d408c109f1f7100a0b;
mem[315] = 144'hf3af00e0f6dffc180139fe7b060cfa8b0902;
mem[316] = 144'hfda9f15a0dc30bc2f67bf57bf4ab0524f4bb;
mem[317] = 144'h085c0735f9300c58f43f011ff6d0fb16ff78;
mem[318] = 144'h01c4fb2b01a4f2ae0221f6900157081dfeb5;
mem[319] = 144'hf2cc02a4fc8903bdfcd90e77f50cf28ff246;
mem[320] = 144'hf8d209d203d6f67b033205d90ef0083109d9;
mem[321] = 144'h0572f9c7097f0d66f10ff2350e420e340b4d;
mem[322] = 144'hfe79fb6fff41faa30de800c5fa22f810f6f7;
mem[323] = 144'hf0740392fd6004a2f187fbdffc1203a0f807;
mem[324] = 144'hfcb8f884f1560d1cf027f41efe68f4f9fc96;
mem[325] = 144'hfabbf77a0acff4570702f3cffa6b0e01fc9e;
mem[326] = 144'hf9180e690d070c9308b9fab80e98fead05eb;
mem[327] = 144'h06740c7dfeb0fd06fd68f598f0d2fb55f8cd;
mem[328] = 144'hfee50c29f343f07bf397fee5048f0805f954;
mem[329] = 144'h0e400ee4f4a4f17c0771045206690d9e0e58;
mem[330] = 144'hf9d30c43fa5100d4f4c7098c08c40fb00e7e;
mem[331] = 144'hfa610efcfc54ffd4f7320e7cf09006e70286;
mem[332] = 144'hfb3cfb920f0e0afd032ffd040624f8ab0be8;
mem[333] = 144'hf60e08aefeb3eff1fe3af6c806daefd60c56;
mem[334] = 144'h04cc0499fb5c0f53005e0ada08dbfe56075e;
mem[335] = 144'h028bf2b8fb84069a0a99f7b1fe91f56cfbd6;
mem[336] = 144'h00cbfb4a0dad0817fd5af6c1f666f3c60346;
mem[337] = 144'hf92df0290326fe3df84b07360d5100b804e7;
mem[338] = 144'hf50b053d095d0ea10b190366f882f70bf90a;
mem[339] = 144'hf961fa30f7d9f1e70a8a042ef2fcf284f007;
mem[340] = 144'hf1a50a320d9901b304e6ffbef717f7fd0fb0;
mem[341] = 144'hf198fe89f3280271f60df06a0cefffbaf4b2;
mem[342] = 144'hff7cfc57f3960cab081d083bf78bf6a1013a;
mem[343] = 144'h086af0d70ce306830b03039105a9f110f72f;
mem[344] = 144'hf37a038c0f05fa3ff8b7fa79fd1bf90cfc35;
mem[345] = 144'hfa9f0d9e0072f9c2f5da02380c69036dfb88;
mem[346] = 144'hf217f4ecfc9e098202830e3ffe170fb90401;
mem[347] = 144'h04dd0e550906f035f8e7fceb0609f236fa35;
mem[348] = 144'h0d46fc05f6250d58fc7ff9b307e4fcfe00d9;
mem[349] = 144'hf7c9f87ff12503ba0f93f61ef6e2f4fc0378;
mem[350] = 144'h02db01730036f2310cbb048af4c902770af8;
mem[351] = 144'hfc2ffffcf5b100b8f396025df86df09c0e14;
mem[352] = 144'h080afaeef71f080303f5fea1faacf025f9d0;
mem[353] = 144'hf91e0c42fb0efc72f4630e0efc20f7c8fa7e;
mem[354] = 144'hfd7dfa12fe9efafbf4610875feb2f7800d3d;
mem[355] = 144'hf7b0f9ae0df10d6e0606008d0f0304a9f2e4;
mem[356] = 144'h0e56f69b080b0b670e920adcfbe2fc99fec8;
mem[357] = 144'hf68afedc0a66fdd9fea9085f04b406600c41;
mem[358] = 144'hf667f8530f31f852f64805b3fbe9065cf435;
mem[359] = 144'hf8a6f76801520537f07d0fc90b2f0cb501c6;
mem[360] = 144'hf43e0edef4ebf6b60541f647f72aff4c0c20;
mem[361] = 144'h0540096efdff0c140b3d01ed0fe9fb5d0027;
mem[362] = 144'hf46e0846055cfde702c2f56908220a95f18c;
mem[363] = 144'h08f3fab800c3f05ff56bff9c0c36000cf478;
mem[364] = 144'hf4e502cc049e0b3a093d0428fc21fa6e0a69;
mem[365] = 144'h075702e1f09a003c0270ff8df10f0857fb5d;
mem[366] = 144'h0b7ff725f3610f6f0ce5f03f02540e0bf4f7;
mem[367] = 144'h097006dafd7c041efb91ffc80cacf3710f33;
mem[368] = 144'hf4e207e1fdaff1d1f5e202e601a10e1fffc8;
mem[369] = 144'hf117091bfa3bf7340ab700960be2f90f00bf;
mem[370] = 144'h03050c3dffc2f2010524033503e809e4f753;
mem[371] = 144'hf665f48709abf57e031204cef5faf5a3030f;
mem[372] = 144'h0c0b04f2f1ee0ea3fff50283fe1afadf0f81;
mem[373] = 144'h00bf0c5cf910f34c0b5f071efd5bfb97fb51;
mem[374] = 144'hf324f68bf69d07dc0c4ef8a705120764fe41;
mem[375] = 144'hf9550e15f4c1f1b707fffaa70891efeffefb;
mem[376] = 144'hfabdfed506350bba0ab409de03c807dc0cea;
mem[377] = 144'h09b7f66807d8f126062ef100fd9a0eedf75f;
mem[378] = 144'hf808f610fd97fb7108c30d1a0d1e089ff370;
mem[379] = 144'h058a07d30365f27cf4fffd65f5c6f27f05cb;
mem[380] = 144'hfa3ff6faf31f0c47ff28001001690ca5f110;
mem[381] = 144'hfaedf5b7fd0f03cc0a310685fa8ff8b2fde5;
mem[382] = 144'hf10cf792fb10f3c50d89f0d00fc9f89e0407;
mem[383] = 144'h0b38fe8c0af4f7acfcabff9e05040c59fc97;
mem[384] = 144'h0e80067d0a85fa59faebf0ce05f50a29fc89;
mem[385] = 144'hfc22fc170f9b0d6cf9eff053026f0d810bfa;
mem[386] = 144'hfa29f975fd9f0399f13d070809720655f7f3;
mem[387] = 144'hfb110afa085ff2cdf6de0be1f51103cef993;
mem[388] = 144'h0a77026e071b09c30358f8d1f1cc0db2fff3;
mem[389] = 144'hf797f88b00cef068f4640b360a85faff027b;
mem[390] = 144'hf9ba041e0d56fcbffddd03a3f9aef266ffbf;
mem[391] = 144'h0e9b04690bdb09610a3dfe2a02480d35f883;
mem[392] = 144'hf2d902cff402fbf1fbb80abe0b51fa440929;
mem[393] = 144'hf27b016c0ea80ec6f23d03dffabaf9a00830;
mem[394] = 144'hf4a7060b02eef6daf7c10c7bf47809b5088c;
mem[395] = 144'hf96e0382fdf4fa69fd91fdfef560fe73f864;
mem[396] = 144'hf66d0447f687f0c8fe9e0387f9d3fceb0b38;
mem[397] = 144'hff12050309d80cd0f913f235f96d06290b33;
mem[398] = 144'h0a63fa3a034ef852f295f4e904fcfd74035a;
mem[399] = 144'h05cf0701f21d08b200f7f500f501f441f327;
mem[400] = 144'hf59a02d5f7c8020d05a3f42f0ba7fe8cf552;
mem[401] = 144'h0666045f06f1049ef67306c8f60101440508;
mem[402] = 144'h0a59f9410c4e01c3f47ffdae01e90c050568;
mem[403] = 144'h00f4f933f1f3f99b011bfa90fffd0eec08c9;
mem[404] = 144'hfe200205f929fd4b06d5fb95fb6afe730f9a;
mem[405] = 144'h02c4f3b5f2fffc5c0365f7bd0f9d0dde0297;
mem[406] = 144'hf640fb2b055905c8fdcdff390dabfca1064a;
mem[407] = 144'hf693fffe07d0f927f33bffdff862fab40dbe;
mem[408] = 144'h0cf5fbf006e1fa380de607ab0c8bf937f9a7;
mem[409] = 144'hf24af71ffe1d00470db00461f57ff7000934;
mem[410] = 144'h0c120ea7f62b0c46008706660a1a0426f9bc;
mem[411] = 144'hffab07740651f61ef7610d590680067506a7;
mem[412] = 144'h0abff6a6fac3f6cff1c30e90fc630464f9b9;
mem[413] = 144'hfcfffd7af9050acef3db0f00f640f596f25e;
mem[414] = 144'h0ec20321055c037f09aeefda06b501750cb9;
mem[415] = 144'h08c10d290fb4f41e0fdff6850057043f04b4;
mem[416] = 144'hfc86f92c0a7cf8be0c750134f3c40fa8058e;
mem[417] = 144'hf3f609aef03efbbc0a1ffa010fb7ffd70e45;
mem[418] = 144'hf3ed0d060bfa0d01f5e904b0f0cb06c004c0;
mem[419] = 144'hf3fa0d150d03057df1c801d70043056a048e;
mem[420] = 144'h0c4dfa110edc034bf2030119fc0f00d90138;
mem[421] = 144'h0a04f790fe720c31046d03adfc20072e0426;
mem[422] = 144'h0b1af454f72ff01305e2f66cf6030d8500e0;
mem[423] = 144'hfc2d03e408a5f3860eb9f1c20d50f73f0f01;
mem[424] = 144'h052309ac0d0e018cf501094c03410b42f086;
mem[425] = 144'hf1d905df0f050d3501b00175fc16fef7f27d;
mem[426] = 144'hf3a7f246fbf5f16d01b9fe71f9f6f4870caf;
mem[427] = 144'h04700107fe1afad10be6f9d9fe34072c0e3f;
mem[428] = 144'hfee3f23c0803f664f9fdfc820e54068a081c;
mem[429] = 144'h011b0f1ffe6ef45a0173fdf6f77efd67f518;
mem[430] = 144'h025f02c9fe63f913f0a0f5450238f3b508fc;
mem[431] = 144'hfc95036000e30480029bff08008104a4fc4b;
mem[432] = 144'h0155fdb4f8d1034fffe40527f49afae30bf6;
mem[433] = 144'hf260f21c04630c510360fa760c8efd1d03c1;
mem[434] = 144'hf807ffae0432f651047af5a6095005100666;
mem[435] = 144'hf629f38904d7f67efdaef0def1a4fa8cf59f;
mem[436] = 144'h0b4bf496f4bb00bcf5d60e00f99cfffcf43e;
mem[437] = 144'hfc50f810f979f93407d3f16dff6c0a4f0329;
mem[438] = 144'h0635f6cbf4b80aaef39202c206aafdcff70d;
mem[439] = 144'h0554ffd3f77f0c16fd4801a70aa9fb87f6ba;
mem[440] = 144'h02a5fd24077bf67f09f00dca052001daf525;
mem[441] = 144'hfbdf0b74ffcf022f00d10b0e06d406490d9c;
mem[442] = 144'h0dca0ce1fc6afa24fa97eff2f8960d080a4b;
mem[443] = 144'hfe4607bc0929f933f91d01c40fc5f820f6b2;
mem[444] = 144'h0e990527f59b0e65f06af3fa0387f2dafb2a;
mem[445] = 144'h0de5fd5df8d1fe1ef1990433ff9d0c560c60;
mem[446] = 144'hf41cfe8601a2f9480cc00fce0e0e0f61f00f;
mem[447] = 144'h07e6f23500190fdd0ff1fcea0a1ef4c905f6;
mem[448] = 144'hf4f8f76dfc21f3cff5b20f80f290f9350fbe;
mem[449] = 144'hf2c30bcdf36e03f20724fe80f08c0462f13a;
mem[450] = 144'h0df4f666f92408f80b3b0be1f8adfdf50a8e;
mem[451] = 144'hffa003720e3b0f0ff616f703fbb8fe6cf8f7;
mem[452] = 144'h04baf412031c03770c18f9100d6209dcfada;
mem[453] = 144'h08f6f259037a05c2f7faf361039dff7b0672;
mem[454] = 144'hfae9032906b9093301b60b82f32ef770ff01;
mem[455] = 144'hfbe00354f420026300eefe470da40258f4f1;
mem[456] = 144'hf4daf85ff731f31206260997fe23fbdff7f7;
mem[457] = 144'h0417fff3f69206e2fa2d097503caf2a7093b;
mem[458] = 144'h0ad7f28f0018f4760c1af15d0a4cf868f61d;
mem[459] = 144'h03e3f13cf67e0924f3adf258fc7f01560874;
mem[460] = 144'hf0350c910483fc12fd280a0a09f7fafaf017;
mem[461] = 144'h0ed1f6ff0f26fab1f0d2faef0515fae00509;
mem[462] = 144'h08ddf87fff6a0a590b26ff56f5c0fc7c09a8;
mem[463] = 144'h011ffe39f74d04fe0287fdb8f96d09e7fb82;
mem[464] = 144'h0d96f946fdcdfaa8f3e4f877015df55afb07;
mem[465] = 144'h03cb0e320b3e099dfa76089dfd5b0675f892;
mem[466] = 144'h04d3f0b7f934fb070b36f7fc0a3701dc0711;
mem[467] = 144'hfcd1f8f00171f135fa6b09160283f0a8f456;
mem[468] = 144'h00270af7fee2f59e09230479ff2209960754;
mem[469] = 144'h06db0548fb3907780187faf1fd02020c06e4;
mem[470] = 144'h0504fdf9f304f8c60ed2079bf9e7f72af163;
mem[471] = 144'h05b1f355090a03edfeccf5c50c48fdf2fe63;
mem[472] = 144'h02c4f80bf6bff8ae0481070cf493f2c3fefc;
mem[473] = 144'h0a8fff2f00220cd507540bf7f97cf0ca0266;
mem[474] = 144'hfec000080a0c0327f5f9f6adf7850f890bf4;
mem[475] = 144'hf919038509f40eb00a4e0e330af00f2e00ab;
mem[476] = 144'hf4080fa4f5b20d5f04dcfb5e01c7064b0da8;
mem[477] = 144'h04c109aaf97e0fc8f8fbf00bf7ea0f62f75f;
mem[478] = 144'h0f44f881f079047df5aafe2201200017f2b7;
mem[479] = 144'h0a07fcf3070cfd880dc20840f0730638f4b9;
mem[480] = 144'hf61efc98f45301f204bdf30ff699f5d801c1;
mem[481] = 144'h03aef40b047e07d3f0bb06de0aa7f76cf1ea;
mem[482] = 144'h0811f555f7d60eddffc9fb6305cf0f78f08e;
mem[483] = 144'h07810023f994ffad0df6f9240fc8009d01fb;
mem[484] = 144'hf26bff21fcf800930e09f12ef5b3f392fd43;
mem[485] = 144'h0fe100a1034b0caa0dd5ff1103c50712fcf4;
mem[486] = 144'hfc28ff2601b30b1b034b0aeb091ef89d0a01;
mem[487] = 144'h0f23f7830c33f387f8ecf3b008510237f7e3;
mem[488] = 144'h040808b506b6fc4f02390419025bfef5fc07;
mem[489] = 144'hfc44f35af16008f3f9a706c105c90082f211;
mem[490] = 144'hf622fb47f2830d7c02d8ff37f698fe75f7a9;
mem[491] = 144'hfe27f32efba4fb90f4c1f3e4fe12fb4dfa0a;
mem[492] = 144'h0d39055d038b07e2f68cf80bf8e2fe6b0ec4;
mem[493] = 144'h092b039609df0f6003df0bdff465ff0f0958;
mem[494] = 144'h027f0faef850f5e3fccf043909ef099d0e75;
mem[495] = 144'hf45601dd08260703f7b8fd2e0ef70766011b;
mem[496] = 144'hfff50df8f9a8fa650ca30b20f73d03cbf15d;
mem[497] = 144'hfaad037ff331feaf0b1b043f04a80dd5057a;
mem[498] = 144'h09dff99b067e0a8d08f5f9b303340e93029a;
mem[499] = 144'hf9910122f2bb047e0b06f1d3fdde0fa1f47b;
mem[500] = 144'hfb97f7660c2bffe5f99b083af98103c90d94;
mem[501] = 144'hf09805b40b1e06f10e5bf28403530527f5ce;
mem[502] = 144'h014b0c4000baf9a804e8006af47e09d7f658;
mem[503] = 144'h054ff071fb1ef77807d3f454034e013af85a;
mem[504] = 144'hf8ee067f09080675f004f0e50f9b0556f101;
mem[505] = 144'h00550aa307970296f6bff559f83b0c16048b;
mem[506] = 144'hf810f741f65bfce8f44ff1840977042c09cd;
mem[507] = 144'hfc5ff80600fa0ba9f89efc09f1410a880ae7;
mem[508] = 144'hf6110dab07fefc4bf52d096709c503390471;
mem[509] = 144'hf191f05df26cfd5b05baf05d0153febe0764;
mem[510] = 144'h09a9049ff9f20268f1e0ff6109700ec9f058;
mem[511] = 144'h0b7d0896f6b40dc8042502bafd800629fe8b;
mem[512] = 144'hf5c30407088200690b63f0b201f104e7fe2b;
mem[513] = 144'h053ef4a8f968fa7c0546f528fd5cf7750496;
mem[514] = 144'hf1850ebf08c20697f88e0ef0fc2cfa980d6f;
mem[515] = 144'h09cff19dfd42fcf2f80b0658063e071f0b28;
mem[516] = 144'hf75f08f4f6f60b0e0b6ef5f60a8208abf205;
mem[517] = 144'h04dfffa00b31042c031f05bd0987f7b9f09e;
mem[518] = 144'hf45ef05ff6c2f4660561fab3f9defe290081;
mem[519] = 144'h063d0a6900fb0f6df1660e5707c2041d0f75;
mem[520] = 144'hf4defdcafcc6fd6e0b20fc64fb65fcea0fab;
mem[521] = 144'hf8be05a1f0250924f4c00d2bf14df350f56a;
mem[522] = 144'h0a3008a608310ec4073a0641f98c05080d7f;
mem[523] = 144'h0cb807edf5cbf6d3fdc00d6bf8dcf2ef02e8;
mem[524] = 144'hfdf401c6f7960e420639fa11f4b9f69dfc7d;
mem[525] = 144'h0591082b0c970b24040cf61ff30a0ac700e7;
mem[526] = 144'hf7b5ff410d6b0a99f2e6f3f9084e022cf740;
mem[527] = 144'h021b005c04050dfaf41508baf03bf838f155;
mem[528] = 144'hfcc40ce9f0de0082fb610d3e089b0ba40f30;
mem[529] = 144'hfb920d0a086400a5f0aa024d07c8f8460d84;
mem[530] = 144'hfd4108fc0a4cf6cf0eeef624f211f4ddf2e0;
mem[531] = 144'h0d36fdd6fbbcf1d0fc0e044cf082fc95f0f4;
mem[532] = 144'h0b8305d0015f02540a2a004e03c3f915fc24;
mem[533] = 144'h00fef8ee0154057d09c900b002dcf987fceb;
mem[534] = 144'h052d026505450648fde3f5cc08800d1a074a;
mem[535] = 144'hf7e2ffaffcb40b3300860183f9820c6501c0;
mem[536] = 144'h00b7fb9b09bc02df080cf53000ba04bff360;
mem[537] = 144'hfc96f26001f607c5f32908a0f7040835f56f;
mem[538] = 144'hfd6d01ee0bf2fd40f82e09a5fbfff196f544;
mem[539] = 144'h0c6af4b808bcf1f40eae0df5fef50fcef35c;
mem[540] = 144'hfa720607f2a8006b0f59f5b20bf5010409c5;
mem[541] = 144'hf699f7d8f7e50ddb0bf601ddf7c10701f2d0;
mem[542] = 144'hf03803faf8b6f4c200ee00d2f315f37b0139;
mem[543] = 144'hf2a3000dffcdf69df7f6fad60edf0ef6fc81;
mem[544] = 144'h05b00a3cfb2506350b07ff7ff3ec0a64f6a9;
mem[545] = 144'h0f5a052bf9ebfe12ffa7f687f22401b7f781;
mem[546] = 144'h071c05700996f0530f85f2ef0ff3fd56019a;
mem[547] = 144'h0854f6f60b2e0406077204aaf4da02e00b17;
mem[548] = 144'h042cf5280e52f5a20a9202f1053af89c0213;
mem[549] = 144'h0e98009c044c0748f9e00067f8bbff520b9c;
mem[550] = 144'hfee0f1fcfe75f666003ff29bf97cfe19f1ac;
mem[551] = 144'h0bc00031f2f80cf0f50df2e10706012c0afa;
mem[552] = 144'hf82f0baef1d0f9c9f341f96efb3d0edf0a68;
mem[553] = 144'h0933f67af7bdf9daf58efaa403990af0fdfd;
mem[554] = 144'hf939f9150c390e6b02ecfeedf096f14dfc0c;
mem[555] = 144'hf383f8ee06c60490094306b7fd6707a10890;
mem[556] = 144'h0804ff440a89f4350481f772f89bfcc5f694;
mem[557] = 144'hfc220289f7eefe44f7a4f995f2280d7df2a8;
mem[558] = 144'h0ddb0b15080008e506c3fd630ae3076004ab;
mem[559] = 144'hffc40c83ff45fd8ef841003a0c8cf8200bd8;
mem[560] = 144'hf1f7f7fc070df5a50c6df6e2f6f7f0f6fdf2;
mem[561] = 144'h0046f28f086b0bbe02700dcefb43f87cfb4c;
mem[562] = 144'hf4730ae7f81ef6b8f2b30633052701be0dc9;
mem[563] = 144'hfab10d630f7cf6dd09070c3e0cc90257f773;
mem[564] = 144'h0768f48404e8f426fdeff7a603b7feea0835;
mem[565] = 144'h06400d98fa1c0cc1f8b50e17fedd0ea50bfe;
mem[566] = 144'hfe08f95bffb1f5fef75bfed10466fd40fd79;
mem[567] = 144'h08d9f73d095605640a460a720cd80f3ffa6e;
mem[568] = 144'hf28c07e6f5d607490c81056df06ef5750e13;
mem[569] = 144'hf335075afe1300110ad70c84f847f2dff69d;
mem[570] = 144'h0c3ef2e50e3ffe86f186fcbc0307f8e004c4;
mem[571] = 144'hf0d4f14d0b14f19a036aff94f6930e98f7e1;
mem[572] = 144'hf62cf583012efcb304770dcd0f5efa0a0912;
mem[573] = 144'h0b49fcd705e9f48cf67bf8a203ac01250034;
mem[574] = 144'hfc5af7c805390599f6b70ebc021d0a94f626;
mem[575] = 144'h0f15f83108e50073f5130ddb0e1aff03f61a;
mem[576] = 144'h0fdefc57fd12f4c1f298ff7f0aaaf7da01ae;
mem[577] = 144'hfb49f25c0d98f03b02f202a90ea4f514fa70;
mem[578] = 144'h043dfd5e096300fcfa52f2e6f755f0c3f631;
mem[579] = 144'h0704061cf1aa0421f05ff540f17b002c0810;
mem[580] = 144'hf5000566f1170508014cff8bf85cfbe10777;
mem[581] = 144'hfef50818f2450da7fd8af433fdd604900998;
mem[582] = 144'h08d4ff5efebdfbb701a0f2c3071402aaf252;
mem[583] = 144'hf478f5a0f7be08c9084fff39f165fc60f74f;
mem[584] = 144'hf175f932f896facffb520c2bfdd9f3e00a7b;
mem[585] = 144'hf4ecf56a09eb0783fa960aebfad0fa360a02;
mem[586] = 144'h0bc400c00978f24bf337031000cef239fef9;
mem[587] = 144'h055a051dfca004a702c7fb590a8a0f6bfe04;
mem[588] = 144'h06dffbd3f2480bac0aac0431041dfbbff39c;
mem[589] = 144'hf8f0f4d80204083efe8ffa91f2760885f353;
mem[590] = 144'h02e7f470ff34fd1d0128f62cf7cd0d8e040f;
mem[591] = 144'hf12a0b370d87016b0661f2f4f9650d0604bc;
mem[592] = 144'hf988f3ed0a3206ad06f0f32ffae8090ff6f3;
mem[593] = 144'h05de0c9f0dab0dc4f8cb028f0de2f823011b;
mem[594] = 144'hf7e5067f041af37cf878f662f2eb0bba00ce;
mem[595] = 144'hf10df3a5fb6efca0f7130555f0eff48cf1ce;
mem[596] = 144'h0e5e0512fc71f6c90d3c0d750be8ff3afc32;
mem[597] = 144'hf97efff3f039fdf4080104c4fb7d05d20185;
mem[598] = 144'hf380f57108af06e102e202d906bcfe1f006f;
mem[599] = 144'hf81b0d77fec50d4cf4db0d14fafbfaa00724;
mem[600] = 144'hf265f8830e680f3cf4d9f220f7f10d4ff525;
mem[601] = 144'hf1a6f98f0ae0012307daf66efec9f55508a1;
mem[602] = 144'h0a2bfafe0c2706f4f6290381f0980426f343;
mem[603] = 144'hf41d005803960479046b0d750a16fb9efa30;
mem[604] = 144'hf7030919ff40f9ea083dfe23f690f169f8a6;
mem[605] = 144'h00e20664f6e007f607e40acc00c008cd0b2b;
mem[606] = 144'hff9cf927faa2ff3905ef0bb20e72fe680133;
mem[607] = 144'h0adf025cf9af02130d2301590043025b0758;
mem[608] = 144'h05a509e2f09302b5f8f6f23af8aafcaef35e;
mem[609] = 144'h0414f63a017bf60ff3e20588fe300b2b0822;
mem[610] = 144'h0aa5ff64f7640b16f6e60354f77a0c63f3df;
mem[611] = 144'h03a2fb6f0fbc093df1e9fc090227f94d066d;
mem[612] = 144'hfcca04850bbbfe400320fb99effdfe050ceb;
mem[613] = 144'hfd3a0c4f046efb56fe9a0adf0cef0ddd05cb;
mem[614] = 144'h05ffffdbfb8efd5909c70ac4050bf24401fc;
mem[615] = 144'h01960e37f90df62c0b26f604f762ffd8f468;
mem[616] = 144'hff1fff26f514fcfe090df42a04e606e7f5ff;
mem[617] = 144'hfe1e0bea0ecd063d0ce7085afa000b0bfec5;
mem[618] = 144'hf135081bf4a1f6520157f44afc1bfae4061f;
mem[619] = 144'hfcd0010ffe9504bb09c602defcaaf8c3f01c;
mem[620] = 144'h03f1f78408d90656fa8307ec00d2f38f0287;
mem[621] = 144'hfc180a340d3c0a9af538fb55ff9908020774;
mem[622] = 144'hf6f8040ef0ff02d50d6d0765035a0a950e21;
mem[623] = 144'h09320319047df2d8fab50bcd0c5a059107df;
mem[624] = 144'h0b260ea80876f4870e4df9750c46f2f3055a;
mem[625] = 144'h0fa7f705f81a0ca6f5c209e9f253f3d70a30;
mem[626] = 144'h0a9a0a30fc020d0c088406af0cdcffd207f4;
mem[627] = 144'hf363f996fd340bed06640610fabf0005f5d4;
mem[628] = 144'h035ef5cafc6d07d8f038f208fba6f827f62d;
mem[629] = 144'hfca90d53ff800e150f8dfaf5fb1b0fdd05ac;
mem[630] = 144'hf1e803e406e9f98c09e8f14cfafafe26f94a;
mem[631] = 144'h004001a0f31806f8f95afdc8f232089402f3;
mem[632] = 144'h0137f5e0fb7dff4f00eb019afcbe052dfb84;
mem[633] = 144'h0f5708ec014705800083010efbb7ff7b0d6a;
mem[634] = 144'h05b9f2550ee807a0012f086bfb0e0210f916;
mem[635] = 144'h05ca02ccf95201a30d54f918f6ad0828f1ec;
mem[636] = 144'h017d088ff1b903580930f89c0967f08fff56;
mem[637] = 144'h0e41f32ff4c9078f063bf0fdf4be03a50e9f;
mem[638] = 144'h0630f67a02ae0c470c13025b07050481f6d7;
mem[639] = 144'hfa8c0119f2fc0784f2a0014efb2402630eba;
mem[640] = 144'hf5efffae083901d8fec8fb510ca9fb3b0664;
mem[641] = 144'h0f3105950bacfea60e01f158fbd008bb0350;
mem[642] = 144'hfe59fdc3fe5cfa6ffba70c4df6e7f680f9e6;
mem[643] = 144'hf187f970fbf208ba0be4f97ff6e5f44e0fbd;
mem[644] = 144'h09720a1207aa054bf8b6036102dff4560c78;
mem[645] = 144'hf328fe6df1640e6f0ad5f1f4010ffd2d09be;
mem[646] = 144'h02740757f4fa0572f6affc4a07bb0cd50b90;
mem[647] = 144'h0f2603ce0273f68d06f705ebfe2b028905bb;
mem[648] = 144'h0b81febefa660443f98f0cb60d190a6d055f;
mem[649] = 144'hf314ff82f85e0846fdadfc46fd2306400853;
mem[650] = 144'h0a8d00fafd500319ff81091ef395f00604ff;
mem[651] = 144'h005b05adf6eaf6400c7402d5f3acff5ff1ae;
mem[652] = 144'hf33cf2210157052efc37ffbc0494fb6c0d77;
mem[653] = 144'hfb40f754facaf62a0164f477f9af0a9a010f;
mem[654] = 144'h085a0507f1b400d90464090b0afffaf4fb81;
mem[655] = 144'h08390b65f4b205db02f8ffb2f524058f0a0a;
mem[656] = 144'h0b5ef055fa3cf91a0dedf3a30b9908c3ff6f;
mem[657] = 144'h083f00f507780c4afb0b0c67f154f0a0003a;
mem[658] = 144'hfc660b78ffcbfee1f4bd030fff220700f5c7;
mem[659] = 144'hf18b01f7f3450656f8d704c10cb3fd01004f;
mem[660] = 144'h05be03a307b7f993f466f5920d5ff884f82b;
mem[661] = 144'hff1afa370176f20dfa14f026f6670848f400;
mem[662] = 144'hfbbf0f7affe4fa7f063c00e508b1ffe80768;
mem[663] = 144'h08ba03d2f01806a9ffe60c05f20805cf0e08;
mem[664] = 144'hf9210d9c0a450895fd12f028fcf9035b0dae;
mem[665] = 144'h09edf215f049044af71ef33b0e92fffa0169;
mem[666] = 144'hf82605a7f507f3fcf48bf0ff007cf2310a86;
mem[667] = 144'h011ffa2e09e10947f56c01b9fe7d0b30f344;
mem[668] = 144'h0480f84cfd69fb5f0d5a04cd07d906240105;
mem[669] = 144'hf6d304c90ac80712f7c5f96ff58af89e0c6f;
mem[670] = 144'hfa90fceef741f3a50af20a59f0a90b25fc77;
mem[671] = 144'h0b5cfacc0aee098af3750e19fe50f16bfbcd;
mem[672] = 144'h06270c3bfb2805cefd7100b500a604b8fadb;
mem[673] = 144'h0be5fd1cf6f3f3aaf79bf2defc8b03930fee;
mem[674] = 144'h0ec5f048014cf017f5470b990d1806640f5f;
mem[675] = 144'hf0d6097902defd76062bfb8105db02fa0138;
mem[676] = 144'hf0000dd4f75a08b806ad0433fea7fb26fd3c;
mem[677] = 144'h08d6fac6faf7faeff5b7f036ffeffe4ff56e;
mem[678] = 144'hfb7dfcddf64a0e570c2a04bf05abf550053a;
mem[679] = 144'hf7c6f958f799076807c0fee70cedf44e094f;
mem[680] = 144'hf02100baf4f3f84f076effcdfd6bf925f4f2;
mem[681] = 144'h041bff2e0002013ffc11f5ed02fff966f6cf;
mem[682] = 144'hf2450854f4d5f2e9fa5d08130c560806038c;
mem[683] = 144'h08400beaf352f294f52700020e83f91ffbb8;
mem[684] = 144'h0dc5f3fef4d4ff200b350aa1f188073bf9b9;
mem[685] = 144'hf8d8069efa7d0209f958fbd20e14fef70bf2;
mem[686] = 144'h048e0b18ffa9f06efe910472f28e05fef544;
mem[687] = 144'h02c7f1c0f47508f40073068ff86ff4d90661;
mem[688] = 144'hf04e0ee6026c04c208a30083fec5f0940ea5;
mem[689] = 144'h0f9bf28f07b2025bfe9e0d6ffeccf8b1fd4f;
mem[690] = 144'hf0060fa4facdf9b50c5f056af5f7fe820694;
mem[691] = 144'h0e57fedaf473046ef45b0d12fba809baf874;
mem[692] = 144'hffdc050d0d5cfb5ff154fb64fd57f7f9efe0;
mem[693] = 144'hfee8f7eff050f01e0b13f928f501054e062f;
mem[694] = 144'h06b90c11f5a6f386f849f344f5b0f5f50eab;
mem[695] = 144'hf2970c8b0f77fde5f623f293fe300f3df45f;
mem[696] = 144'h012c029500abf589fbdffe8ff478f14d0d9e;
mem[697] = 144'hff750356f7a203530fb3f169fe1c03dd0196;
mem[698] = 144'h02fcfd5c01640538f101fc280ee3f15ff1d6;
mem[699] = 144'h0afcf00bf2c3f55af0d8fe9d07e9f4bbefc8;
mem[700] = 144'h001efbe40f510179fc9d09d6f728f7fc013a;
mem[701] = 144'h0673f91fff04fbe50a13f66a0a6bfab301c8;
mem[702] = 144'h0427083e099efe28f99100880a160c9cfee4;
mem[703] = 144'h03eaf8e00e090171f23bf7530ef4f0d80951;
mem[704] = 144'h0f8a03c803fff3790705f4000145f49c081c;
mem[705] = 144'h0aa4ff4dfd21ff78fe680d9c0365f09bfb40;
mem[706] = 144'hfcaef8a1f927ff520e0d08f5fe44f5470a37;
mem[707] = 144'h00b50924fbe5f25dfbe2fc4efcbffee4fc0b;
mem[708] = 144'h0f77f7d1f581f2e2fdf9061c04e1f06f0177;
mem[709] = 144'hfa29f75b045dfc650b39f6ca00a6f2d2faf8;
mem[710] = 144'h062cf5e205780d000ae1082bf99900b10c2f;
mem[711] = 144'h09a1f067079c0b6c09ba05b600d20a9e07fd;
mem[712] = 144'h03bc0b9cfc020f07fa670b44ffeb0b6509cb;
mem[713] = 144'hfec8ff93fdae095ff8fbfe7af8ab0423f38c;
mem[714] = 144'hf0faf7b7f5c9fd89f1fefd39074c004801ee;
mem[715] = 144'h0d0c0a1904130213fa9300460f9bf03407a1;
mem[716] = 144'hfe7e0a000b44faf7fcbbff2df10b0a72efb8;
mem[717] = 144'hfe29f86f03ca0d1bfc5a0dd20456001ffe0e;
mem[718] = 144'hf2ca0f90f3bd0bf0f70b02ff0509f35bfd7c;
mem[719] = 144'hf54bfc97fb7aff390a65f216fa8e0a6507bd;
mem[720] = 144'hf89efe5df042fad301f709dd09c207030723;
mem[721] = 144'h0e37fbd7f97501d2f744f82afb37fcd5f5dc;
mem[722] = 144'hff9bf1120686f8650082012e03bc096605df;
mem[723] = 144'h0833fd530df6fc2f0ab305b2f68f05920060;
mem[724] = 144'hf039f17e0a91074405c5f1c20874fe5efb0a;
mem[725] = 144'hfc64fb9701a2035af399f9b106de05f60438;
mem[726] = 144'h0970053a0c870d8109c2fc90fa0b0d270daf;
mem[727] = 144'h0683f577f2df08d20b36f2ea0f17f130fd06;
mem[728] = 144'hfbedfe120e1209aef55404a8fc59f1fdf57c;
mem[729] = 144'h01380a71f06b03b0f4340ded0834089b0e64;
mem[730] = 144'h012ff62bf989f825f130fbb300f6f59e0e8b;
mem[731] = 144'hffb7030908a4f86d07d8ff0af073033ffdb2;
mem[732] = 144'hf550f8910afd006ef4db0786f35100190466;
mem[733] = 144'h0767fa92fbfcf763fa120ed105d10cfbfc62;
mem[734] = 144'hf8be0b0b041a0c18066ef9f703fe064c00f2;
mem[735] = 144'h021e0ee30676fc310f5103dd0e77052ff949;
mem[736] = 144'h0a5201420addfd5a05f50650f8d9fa990440;
mem[737] = 144'hfb3af818f2ec0fd5f1fcfdee09650690061b;
mem[738] = 144'h03c0f4b80db405a9f05ff01403010c5f0609;
mem[739] = 144'h02c607910642fdee06380809f79908320062;
mem[740] = 144'hf14cf12dfd2506ed01a7fa75fc260cf204a8;
mem[741] = 144'h0695f8e0fd14f476081b02e6f980f8e60a58;
mem[742] = 144'h0291ff810334f03efbb4f1200fcbf0ee0695;
mem[743] = 144'h0d800136f1fef5fbf4d3f1cc0977f212fb66;
mem[744] = 144'hfed7fa2e0e40fa33fbd4f9d7f9a3ff660242;
mem[745] = 144'hfb8ef15e033df1a7002d0106fccd045f083d;
mem[746] = 144'hf701f9fc0724fc6d01d0fa230ff70851fad4;
mem[747] = 144'h0bb90f500e29f927f0e801f900e505b0f72d;
mem[748] = 144'h05d0f28f0ae20e12f17e0507fc43fee105d8;
mem[749] = 144'hf292fef307a30d9f00520c100450013d0f08;
mem[750] = 144'hf3e20d0801a8f19505c90b76f90af68900a2;
mem[751] = 144'hf436f3f9fe2c07cafbb7f792052b015bfd86;
mem[752] = 144'h0658fbc8f05a0c5ffad9f424f434fcbcfe4e;
mem[753] = 144'h010305c109080ca3002601fd0fb10db20853;
mem[754] = 144'hf23dff5803030d27fd6af65b054ef48f00fc;
mem[755] = 144'h07a5fb70f7c6fd05063cf6610c4cf5d3ff00;
mem[756] = 144'hf34f06fc08a6f298f5b1039cfe8705060dd4;
mem[757] = 144'h0cb70f8a09c0fcfcf46f020902f6f780f83f;
mem[758] = 144'hfe8fff09f84ff113076cf2000925f53df2aa;
mem[759] = 144'hfce1f35e095ffdb7063f0f9b00c8f2b10cc6;
mem[760] = 144'h0a2b082a0fcefaa402dbf1d808e20449f22a;
mem[761] = 144'h05dbf9b0f8bffaf6077af0d6fb9c063ffdb1;
mem[762] = 144'h059afcc00ec0f9e6010afe63fb1103100a50;
mem[763] = 144'hf47df9180caff91bfb24052dff310fb9053d;
mem[764] = 144'hfc42f1320995f79e00d20ac1f0d4f58cfdb5;
mem[765] = 144'h0aedf88c0cfd02cc02e4053ff302fc51ffec;
mem[766] = 144'h09a1ff720c3e08b2f0c9f7eb0cbb0907fb09;
mem[767] = 144'h0bc907590479f0cc00ebff6c0d23f2200833;
mem[768] = 144'h09e20c5ff579f9870549fd35083e0769ff66;
mem[769] = 144'hfc06f4eb0bfe013a080affbc0cadf1e9fc74;
mem[770] = 144'hf4900c7102fa0241f3e8fe0af8900e11f60b;
mem[771] = 144'hfa380e6407bff8c20b4e05b40d7a03d4f4ee;
mem[772] = 144'h034ff7cafae10791f2bc0f73049af49602ce;
mem[773] = 144'h0829ffbff510f26a036bf6f90b02f84b0bb9;
mem[774] = 144'hf60bfc5002a301010234f051066af4fcf823;
mem[775] = 144'hf82af13ff024f27003f4f77bfa39fa3ffea0;
mem[776] = 144'hf2a90adefc11f69afafef3f7f3fd06fc0f20;
mem[777] = 144'h0de6f0420d1300eafa1f0407fd46f538007d;
mem[778] = 144'hf09bfab10435facd02c6f045fbb00caaf275;
mem[779] = 144'hf84f02180285fb1608c9fed20e6709c80793;
mem[780] = 144'h0241fc43fee8065af2cb024ef92ff4d9f9d7;
mem[781] = 144'hf92302bc0f670025f629f0a6f44f0f26ffa1;
mem[782] = 144'h0585ff3d0fb00aca04fa02f701e70195fb7f;
mem[783] = 144'hf8e30f4d0624f85e00e2f167f40cfd1d0761;
mem[784] = 144'hf8ea0e98f357016dfa4b05fbf3befcf6f2a8;
mem[785] = 144'h04370d90f37af32b008c0566f40bf24bf0cf;
mem[786] = 144'h04eff911079af8780e7501ddfd90f002ffc6;
mem[787] = 144'h0b230801fa73f767f96d094f090308a3f6e2;
mem[788] = 144'hf17af4a90c85f2aef5fafe8c0786f845f856;
mem[789] = 144'hf457061a080d039e0959fc7f0cd90f040e6d;
mem[790] = 144'hf54cf4b6ff43079afa24026d0ab1ffa0fb21;
mem[791] = 144'h07adfa43f6d6f584f00309fe0ad2f52af550;
mem[792] = 144'hf227027cfc2605c8f8b80e21013cfb44f772;
mem[793] = 144'hffb10a6f0b6ffab9f20604df01570ed7f8bf;
mem[794] = 144'h0b13f827f6b800a2f7e3fcaaf05a0a480201;
mem[795] = 144'h062ff2060430f6abff98fbe30461f95ef658;
mem[796] = 144'hf7180676ffbb02ca0abff1df0cbefefcff65;
mem[797] = 144'hf0340ca10b9dfce0067ef8e8fa3bf0340b27;
mem[798] = 144'hf5fefb99f11a08200c0ef9600f67f6170533;
mem[799] = 144'hf59f0389f69708caf75b0c02fa13057b020b;
mem[800] = 144'hf2b70b33ff70fcd3f31cffa2089f099dffe6;
mem[801] = 144'h0ff103ddf942fda2fadc0668fe91f798ff8f;
mem[802] = 144'hf6f608e9fbb10d7bf871fc1e0994fdf201ac;
mem[803] = 144'hffa8f068fbad077104b70724f7b8fd3f047c;
mem[804] = 144'hfd71f1410b560c88fbccf81b044009220cc1;
mem[805] = 144'hf3c0f4bdff5dfa67f68bfa9608f30917fe59;
mem[806] = 144'h0bdc09eb0b8e05f8fa4c0842fb84fbf60c75;
mem[807] = 144'hfce10d3cf8850277ffa0f45af1f0f178faca;
mem[808] = 144'h0a0f05190530f60ff7ca0bbd0b3f069c0c2b;
mem[809] = 144'h02600d35fd7b022d0b8302e1077f04f2efe2;
mem[810] = 144'hf6ca0293f3fdf72007dc003bf02905290e25;
mem[811] = 144'h0fabf9d1f771f9d6f2caf5350d0afbaff3cf;
mem[812] = 144'h00c50af6f54c0084f4a3092802fdf9580cd6;
mem[813] = 144'h08000c490cba05230dd8f117f711f78403e6;
mem[814] = 144'hf1cb0d31fd3bfd200d6ff900fed0f37e0eb8;
mem[815] = 144'hfd78f66cf498f8620d63078e07850dbbf858;
mem[816] = 144'hf0b409effb72072ef1c504060d41f81df6a6;
mem[817] = 144'h01cd090d077ef5500d6a0cf5f0a0f3b1f17e;
mem[818] = 144'hf3cff573fe81f20e0c9804b30dd5f05b0a81;
mem[819] = 144'hf3ac082affc40c24f98ef59b02acfe0c0365;
mem[820] = 144'hfb6309e1f4380c6b0dcbf130090d0746f08d;
mem[821] = 144'hf30dfe2ffd73f2b9f10607def6ff0698fa70;
mem[822] = 144'hfdb1f38705a0017bfcb5f2c90a8c08ac0701;
mem[823] = 144'h0141068d0683fa77fd410937f6910f69f19c;
mem[824] = 144'hf808fe93f407f8df0b6afd7afbdc00f804d1;
mem[825] = 144'hf9670e4df6fbf775051500370f54f7890a3a;
mem[826] = 144'h086804caf12c0fdd08c40a6df6ab03e30001;
mem[827] = 144'hf127f1e9fec6f6a7f3400d7dfba2fa300fc3;
mem[828] = 144'hf5e109fef43bf915fb94f6f8f1cf0260f34a;
mem[829] = 144'hfa79f96cf214f7df0c090fff0bc6f5230f95;
mem[830] = 144'h0c4ef1ebfc16f66f087df308095201b7fd39;
mem[831] = 144'h018dfe33fc9af15af6de0b510c86fb6c060e;
mem[832] = 144'hf67202d2fbc107d7fe7709460f30f89c01f8;
mem[833] = 144'hf157f217fa680bbaf246003d0f3df25afec6;
mem[834] = 144'hf1600766004c04010ca302bdfeeef781f677;
mem[835] = 144'h09fe0d2cf66a08b80e3af34df675ffa4f5d3;
mem[836] = 144'h06530ae705d50238064a0212f1190a56f74b;
mem[837] = 144'hf8b7f4f205b507fe0984fb9f04310f41f4f8;
mem[838] = 144'hfd100a0b036ffa5ef33df203087af480f859;
mem[839] = 144'hf4fa045f09b70a5af1a80131f8fc0623f2f6;
mem[840] = 144'hf760f3cbfd48044500f6f131fb30f5ecfcc9;
mem[841] = 144'h04ccfa08011cf4f5f4a1f22b07acf6bc099a;
mem[842] = 144'hf797ff14fb2bf1ee015bf7ea084d0f81fb02;
mem[843] = 144'hf2e0f6a5fa58fc330697f64b0fa6f5a0f586;
mem[844] = 144'hfafff0c80b1805aef8980dff062e0ea90050;
mem[845] = 144'hf012f72e0a62fb150b520790f6f9006df46e;
mem[846] = 144'hf29d0fc5fc27fba8f7b6f72efad902810c15;
mem[847] = 144'h0b94f1aef0bffbddfc12f044033dfe20f69b;
mem[848] = 144'hfa73f721ff86f12004510e3101ebf455f794;
mem[849] = 144'h08e4f51dfca50dd7f160f964060cf5bc072c;
mem[850] = 144'hf538f7c80d870e3008b00863f9bf069300c9;
mem[851] = 144'h0544fb1af92af12108fa0a26f402f6e60bb0;
mem[852] = 144'hfb9df758f4c90b1af552f176f33a0df606f0;
mem[853] = 144'hf182fca20f9b07acf109fd6706be05f709c5;
mem[854] = 144'hffd30a150c1c0272f8a9047a04a00560f414;
mem[855] = 144'h0edaf28c04ea078a01fff7860755068bf509;
mem[856] = 144'hfbb3ff29f3d7f30f04bf08e40ecaf3acfd20;
mem[857] = 144'h0c7a08ec05b208240491f4990f280f2706ec;
mem[858] = 144'hf228f96cf5b6fb1c0aa3f03209400259fffd;
mem[859] = 144'hf0c704070a070307f2e5f8b6035afa41f6a5;
mem[860] = 144'h0f410432ff23043efa31f110f4380dc5f328;
mem[861] = 144'hf5060c55f62e0365f5dafd1af73f0919f003;
mem[862] = 144'hf91efc2c0282fac00fe00e87f6d2f8a6f810;
mem[863] = 144'hfde403e4f729015e08830725f54907e10b01;
mem[864] = 144'hfdc1f6cdfd4403aef0de09a9f8960234fc44;
mem[865] = 144'hf47c0d5500e6084df1af0155f4460bd20441;
mem[866] = 144'h005af29efe6c00860d15f596fe0f063609d9;
mem[867] = 144'hfc37f246f95c01bc0a660f5c06010aa700e3;
mem[868] = 144'hfa6207eefd21f40d08c00e02f155f617f330;
mem[869] = 144'hf54a03180f75f76007ba0249f01af68a09d6;
mem[870] = 144'h01c1f89509b70cb7f0fa0cf4f0fd0267084b;
mem[871] = 144'h0219f75fff05f03d0bbdfd170240f7820437;
mem[872] = 144'hf06101a20045f294f871fa48f9f004a4f4de;
mem[873] = 144'h094a048f0723f4b2f6330c19f489076ef103;
mem[874] = 144'hfdc403eef0d8f90af6bdf8edfaf0ffad0100;
mem[875] = 144'h060607f5fb25043105a9f7a9f54ff66300ed;
mem[876] = 144'hfd270e010d7ef96e02f70c500471077e0cf6;
mem[877] = 144'h0c5901a20d5f08bdf6effd3f0221fab00494;
mem[878] = 144'h0b75fc38028f0e8efa2af296025709d90f76;
mem[879] = 144'hf446068cf1930ac0045706f8fca604b6ffbc;
mem[880] = 144'h030ffa1ffa6d0facfb85f44103c502ed0984;
mem[881] = 144'hf6a8083900d3fe06f9780b36f86d0b3af5e3;
mem[882] = 144'h0b970b2c04380e6ef051ffe2f9a5f865fb33;
mem[883] = 144'h06e60b57fdaf02bc078807fd0cfb00040f19;
mem[884] = 144'h05a7f9050199f68cfd38fe86f50700dc06f1;
mem[885] = 144'h0ee80ad00fb7f9d9faa302970330003c05cd;
mem[886] = 144'hfd6ff2e703090c5f04f8fd1c0fce0a0009a7;
mem[887] = 144'hf3fafa0f083808610e57f51003c808e8078f;
mem[888] = 144'hfc35006a0cc4078f0c6f03fdf704f40ff096;
mem[889] = 144'hf04204a2fbb3fe460c94ffa1f6b8fee3046d;
mem[890] = 144'h02cf0c4c0505fdb2fd6ff15df1a804fc0d81;
mem[891] = 144'h0345fff4f8f4f6d0f53208e6f35b00b3f20e;
mem[892] = 144'h05aa0027f3c90589fa9ef64a062a09840d11;
mem[893] = 144'h052ffbd9fe0ffd98f2bd0b010567f8f1f5fd;
mem[894] = 144'hf18903980f83f206011bf1d1f119041704d8;
mem[895] = 144'h000d0f28fc190d0f09ac0e0d0b6afa09f266;
mem[896] = 144'hf1f20761fd3d0f24f5610ba3fec7f8e4efe7;
mem[897] = 144'hfb2af8cc087e0aaffdd40f020e750b31f984;
mem[898] = 144'h087905e7fe8ef8a50e82fc28f8a9fa44015e;
mem[899] = 144'hfd5ef2fbff42f7da09600d1407f8f340f918;
mem[900] = 144'h02aafad101a8f19506ac0bd40ab6f8faf7aa;
mem[901] = 144'hf59e0ce50062f4ecfd19f0d10e06feddf6eb;
mem[902] = 144'h09380199f5b1f9970cf208f508ad0334f846;
mem[903] = 144'h00e3fce802aaf4dc009bfe16f80d095308b0;
mem[904] = 144'h09cf017f0631fa8a0ede06a60de408d0f265;
mem[905] = 144'h0450f452055ff9380f280344088b04bc01d7;
mem[906] = 144'h0f0e0be7ff7bfafff3bbf23cf62309aef78a;
mem[907] = 144'hf034f1e602c9f5f3095501f20faef029f9e1;
mem[908] = 144'hf3bff54204510c28f6480fad0948f606f3f4;
mem[909] = 144'hf6e7fbd00235fbc6fc7df696f06ff78dfc36;
mem[910] = 144'h09e8f97808390a950f730e31fb2f05e7f6e1;
mem[911] = 144'h0890083006e303310035fc3c0b53f90afe38;
mem[912] = 144'h0ab2fec70618fcc0f6cf00a1f414fbd3fbe1;
mem[913] = 144'hfa630d300e2fffe8f88ff55303fc0180fb5b;
mem[914] = 144'hf41e0e6e019d009cf25d0f09f435f2bd06b6;
mem[915] = 144'hf1b2015f0db1fc87fcdb03520a19fb6c0e59;
mem[916] = 144'hf7a2fa7808850625fa9e0da101acfcd5fd33;
mem[917] = 144'hfea9f45804e4f111f5eff2adf29efeaefa10;
mem[918] = 144'hfd260a560d91f83dfbcbfff9fa3e07220982;
mem[919] = 144'hf75bf314076b025c08c2fd6df52df4f8003b;
mem[920] = 144'h08aff94f00b80388fdbb0c5e04f7f5a2f4a6;
mem[921] = 144'hf1f20cd0f604f00b0137fff10dd1f6edefe5;
mem[922] = 144'h05c40a6e0a660a4605ecf2a90276f4760493;
mem[923] = 144'hf35b0a78f6ce0a98f6750e55f858f46bff81;
mem[924] = 144'hfff40405f48d0cf3ffa1fb3c0470ff66f6d2;
mem[925] = 144'h03470cd3f4d1f6fc0818f68b0e540e700d2e;
mem[926] = 144'hf95f0458f907fe46f72d067b063b0d88f6af;
mem[927] = 144'hfe23081506a9f22ff222037604af0d3ef2e5;
mem[928] = 144'hfc76f82ff45df13c0a4ef4adfd1ffc6ff3b4;
mem[929] = 144'h026cf0f1f27a0661fe69f172025cfd95fc6f;
mem[930] = 144'hf20f0f7cf14e0cf3f9110df1f51ff11ef676;
mem[931] = 144'h02b50d250a8609caf422fe8ff7310a3f035a;
mem[932] = 144'hfbfbf214078ff96201a205cff57df7a9f942;
mem[933] = 144'h06ec01bd09df01a60e1bfffcf6fc0e1bf173;
mem[934] = 144'hf6d305a204f00543f83ef85df12a07c0fda4;
mem[935] = 144'h0b6406e303a10f46f12efa0af76efc21f0a7;
mem[936] = 144'hfc4cfc3203c7fef90bfafdd3fcc201820f2e;
mem[937] = 144'hfd290a37f84d0dd2f85ffa5d0a670ea80fb2;
mem[938] = 144'hfcc10920f1defff70c6b03cb0d5ef35402a1;
mem[939] = 144'h0c73fae309dd085504c3fbe00a220239fbed;
mem[940] = 144'h081906280f9b0c7ffaaf0ffb0e1408d107c4;
mem[941] = 144'h07a7f633fc27f8880a640c470a060caff928;
mem[942] = 144'hfef30acbf7e1f49ffa74f74ff0dcf698f3c0;
mem[943] = 144'h0dae07750650f08afcfc0f56febf05c1f3be;
mem[944] = 144'h08b4fb6b0cf2fa16fef5f02805f807ab0e31;
mem[945] = 144'hfbdb01640c08f0d80e3ef59ff3d50c800e3a;
mem[946] = 144'h054800e0096ff6baff620c57ff960815045d;
mem[947] = 144'hf953009bf928f985f4eaf169fc24f3d0089e;
mem[948] = 144'hf651f2550d0b07ee0fe3fb690dcefb70f4cd;
mem[949] = 144'hff82fc25f6fc0535f4090d260d5302c1f50e;
mem[950] = 144'h0499f7f6062cf99e0bc9fc05fe8c03950c36;
mem[951] = 144'h0d320a63f8d6f008f4240de7f2adfba902ed;
mem[952] = 144'h0a4afc18f38407b60b260e97fcba03b7f51f;
mem[953] = 144'h0daaf7620377f2d5fe2a0444f74df7fc0da3;
mem[954] = 144'hf18200b8fa94fac1f4a90574fb9c0f2bf79e;
mem[955] = 144'hf8d6f593f1c4f960fc74f182f794f102020b;
mem[956] = 144'hf8820ee7f7a9f0490b3df4e70bdf07b8f639;
mem[957] = 144'h0e56f8bf0574024d0da7f56af4760e8a085f;
mem[958] = 144'hf3210d2a0eec0683f1ddf273077bfd3ff51f;
mem[959] = 144'hfc2907b201fbfd70f9cffd0cf1f0f1cd0c02;
mem[960] = 144'hf14df82a09b805a90082fa940c57fd8f0782;
mem[961] = 144'h0e9b07c40835fcc309890c430577f27cfd50;
mem[962] = 144'hff650cf0056b0a650efffe21f2bdfa5cefe8;
mem[963] = 144'hfd0ef1a00ea0ffa10a1b0327fd5b04b8f203;
mem[964] = 144'hf841ffd5fed6011c055909a70155f542f9e9;
mem[965] = 144'h01eff99505490f6ffeddf7c3f667f50ffc67;
mem[966] = 144'h0dbcf89b09ac044007c3ff1c024af7db08d8;
mem[967] = 144'h02a80678f3c2fd9df0cdf7cd0b500962faa5;
mem[968] = 144'hff56f93ff42e03f7f52b016cffa206260724;
mem[969] = 144'hf118f49a0535fea5f011f10501950fb607e8;
mem[970] = 144'h0461f03afcf90c76fe1ef9adf7e10a54f5be;
mem[971] = 144'h0ed1fb21f364f2c8ff3903e70a1201a4fc13;
mem[972] = 144'hf5e6094e0b13074903a305b90794f1a10282;
mem[973] = 144'hfae304ae0d180a91ff91f8cdf57a07e7fbc7;
mem[974] = 144'h0690fcbbf0d80886099e0a9ffa26fde3fbb8;
mem[975] = 144'hf0b6f391f6170bb50c8c0ec304c402be0f89;
mem[976] = 144'hf1e7f826f88f044f0de40da3f13c0c93f198;
mem[977] = 144'h0ee4ff8e081e010d07f90474019203a50966;
mem[978] = 144'hffdaff3ff669f4610213080c0da000b2006b;
mem[979] = 144'h02c1fe1b07230900f0fa09010df1079202e8;
mem[980] = 144'h0b1dfc08fcd3fa7e0c7202700a91f0140445;
mem[981] = 144'h082c07fa00780ca60b3e04e4f9b20ee40c90;
mem[982] = 144'hf667f8b3fc0901eef887070500d6f489f879;
mem[983] = 144'hfae907d2ff41fe460a040ff00c23fb8808fa;
mem[984] = 144'hf798f042fd33f99bf09705f4fa9e0b90f70c;
mem[985] = 144'h08ef0987015a063afc4ff1ee03dd0afb06a3;
mem[986] = 144'hf2fdfca1f9e5ff880fb40d84f4480715f17e;
mem[987] = 144'h06d2f458f47ff27b0157fee603bd0b92fc8f;
mem[988] = 144'h0e33fd3808f009e00f230776fccb06a8f3cc;
mem[989] = 144'h09840092f55efec7f2f1fbe4fdeffee2f385;
mem[990] = 144'hf6edfc7dfe4f0f06013ff7d5f917f5eff01a;
mem[991] = 144'h040df3e708b604e0fcb9f8fa020af63f0628;
mem[992] = 144'hf3ebf1bc0cc90410063306920fc4fff902e7;
mem[993] = 144'hfd7cfcb605dff8c1fcecf5cf00e7fb8afe37;
mem[994] = 144'hfa050c52f042fdc6f8870d11f4a00e580205;
mem[995] = 144'hfa1605ec0b71fe6201500a27f35d06840c90;
mem[996] = 144'hfda1fd3f0df90d79fb7405b2fa1dfcd6f07f;
mem[997] = 144'h0ed50f16f76af44bf7adf213058d0339050d;
mem[998] = 144'h09480701f7b9f318fba00254f802ff5af674;
mem[999] = 144'h0fc3077bffc7f1f4fa4df1cb060801b00c4b;
mem[1000] = 144'h08a1f74f066c0d72fcd000520ea1018af7e4;
mem[1001] = 144'h06350ceffc67fc8d01760c9c0eb0028e0038;
mem[1002] = 144'hfa1e0c1a01b60eb201bef0590c21f598009c;
mem[1003] = 144'h0893f18e053004ca04e507d9f9c4060bf0f4;
mem[1004] = 144'h0a23086f0c4ef6b2fbf402b4fbf4f131faf9;
mem[1005] = 144'hf6030bd00cdbfab9f8dbf533f240efe6f545;
mem[1006] = 144'hf367f34d05e20f09f6f5f31cf295078a0a26;
mem[1007] = 144'h0402facefdd7095a0666f5aaf4c4f2260857;
mem[1008] = 144'hf647046d0266f316029af91d0ec80ce40950;
mem[1009] = 144'hfbf8f180f2fdf6980b44049f065a0654fae9;
mem[1010] = 144'hfa28f0b208380be6f40cfbbef4fb0532f011;
mem[1011] = 144'hf495f85d00b20a900a46f72200d6f35e004c;
mem[1012] = 144'h050003d4f30f0a82fde302a3f768f8f203f9;
mem[1013] = 144'hfc61fb2efde4f2bdfd97f04bf6bd0893fa4e;
mem[1014] = 144'hfc4907e0fa7cfbfe088ffef609b1fc22fbd3;
mem[1015] = 144'h0592f02df71eff7b0ce50b6af757fcd3fd72;
mem[1016] = 144'hfd46f5b306abff82fac3f1c80bd90d40ffc7;
mem[1017] = 144'hefe105580d130c650c5cfc280e6208a1f11d;
mem[1018] = 144'h0335f059fe7306c40083f569ff38f21504e0;
mem[1019] = 144'hff97001af389fe9ff60d0c9df0860f470b5c;
mem[1020] = 144'hfa92fba00ac4f4ab09ddf6d1f9fef5fcf467;
mem[1021] = 144'h02a3ff9d03d5079cf098f5020c8ef9d6f904;
mem[1022] = 144'hf087fee2fe35f01e0ed8f5eff66ef820fe7c;
mem[1023] = 144'h0ddc0297f87b04b0f1a5f5770e3401880197;
mem[1024] = 144'hfa020c42f65bf6ac0f75f33c064ceff3f3ac;
mem[1025] = 144'h03d9fa2af0ffff5801f6f7e5f718054d0e4c;
mem[1026] = 144'h0d03f41e0228068af4e1f3b706d0ff190c90;
mem[1027] = 144'h0fa10c9ff1af05a40e2e077103dc0eac010b;
mem[1028] = 144'h00f2053a01e100bc07750d170671f5acf667;
mem[1029] = 144'h04c7001a03f9fb5f0fc90070fe79028b0a5c;
mem[1030] = 144'hfffffb400f4f021c0b03f8470821f17d0992;
mem[1031] = 144'hf59e029d0291f2cf0d88029703980eee1004;
mem[1032] = 144'hf0d3082c038df38007f7fa13fffdf20cf029;
mem[1033] = 144'hff74faf1f8950399f84ff41ff667f8ec083d;
mem[1034] = 144'hfccaf37908200c3f08e6097efad2f2aefa96;
mem[1035] = 144'h0f43095ef2470938f9e40aaf041bfb4bf2bb;
mem[1036] = 144'h0bea0eccf6400e99f42ff8f2f684000af5cc;
mem[1037] = 144'h0c9c0414fd1500c5f1b00177f73cf4cff921;
mem[1038] = 144'hf768035105fc07edf5ad0771fc300cd0f633;
mem[1039] = 144'hf24903bdfb62063cf292f8e9073ffb190933;
mem[1040] = 144'h073108660568083b0970fa8d0505f7b1f4c1;
mem[1041] = 144'hf6590d40f881f7f505e103520b220fd8f5c4;
mem[1042] = 144'hfe64079804eaffadf89500ac056f04940a90;
mem[1043] = 144'hf36dfeb10ea1f2bbfeb8059cf8e8fd700988;
mem[1044] = 144'h0df90452f9f0f3ec0fd30cba008f0290fca5;
mem[1045] = 144'hf18c094f05050b020d9204dc00670600f790;
mem[1046] = 144'h0d160e58f79df18b055f04720686f0fff7b9;
mem[1047] = 144'hf7740638f84707350e1202c4f9cb06320a65;
mem[1048] = 144'hfb85095908350a0ff409fadff3420eaef136;
mem[1049] = 144'hf7d70bd8f2ae0f1a06fc0960f942f7d5f768;
mem[1050] = 144'h0de5f61905fa02b30c4d0b42fa34091ef522;
mem[1051] = 144'hf6c5f7cbf3f4077bf699fa9f0f3dfdf70323;
mem[1052] = 144'h0795012d0df70991f4e5fee107fef368f203;
mem[1053] = 144'h0da0fe0ef4d7ff29fbaaeffd05960f600de3;
mem[1054] = 144'hffd3ff38f4bdf61a083702e7fd10fd8c0968;
mem[1055] = 144'hfd42f4870bd2f295f3def33efac2016ef27e;
mem[1056] = 144'h018d0c3b0aae00740b110279029a0812f852;
mem[1057] = 144'h09d102a1020d04ed0cb0fdd5ffecf6770651;
mem[1058] = 144'h07eefc83044f0381fdc5fae7fb4e054208c1;
mem[1059] = 144'hfab2f75f05660f4df2220eeff65301ec04e8;
mem[1060] = 144'hfaabfadd0e3bf2f4ff40fe9af9230716fee8;
mem[1061] = 144'h0c5c05d704c2066bf125fc65fd680a510cf6;
mem[1062] = 144'hfcd50e68fc83ff36f8d3f1370a2c043208dd;
mem[1063] = 144'h0778f02ef199fa71fe56fc99fe4c081e040c;
mem[1064] = 144'hfdb8f9f202a20cbf0e8a022d01fd0b9c02a2;
mem[1065] = 144'h03360238f50b01f3f17c09e6022cf248ff66;
mem[1066] = 144'h0ecf047e06ecfd3bf34609ef069cf9b1f53a;
mem[1067] = 144'h0fb0f0e6ff77f7c9f144f95c045b0873f31d;
mem[1068] = 144'hf477fb41f673f6b5081e04780e4a00c7f933;
mem[1069] = 144'h03790a760e0bff7ff037f54c0a650c4c003f;
mem[1070] = 144'h06590c5bf9edfa210c3607a3f031f649fac4;
mem[1071] = 144'h0a4aff05f62f07880f9df79cf3dcf48ff6b6;
mem[1072] = 144'hfddc0e43f76cf97302ed089a0f66fcf90834;
mem[1073] = 144'h07bbff200cb007380c94044d035fff800910;
mem[1074] = 144'hf5edfc940776f27afca80b2ef2e5f75d0935;
mem[1075] = 144'hf136f645f218022000b7fd2bfd11f329fed1;
mem[1076] = 144'hfb8c07d503ce0588fa9cf5d4f0e20713098c;
mem[1077] = 144'h0c6cf8500d4cf51a0171fc29ffb2f701f94a;
mem[1078] = 144'h04730325f0d7f0bef6dff1f0faa7f9e1f8e9;
mem[1079] = 144'h01c40097f8e0fe88f622ff88f53af482091b;
mem[1080] = 144'hffb7fc5efc700432f67df718fc32f1820c13;
mem[1081] = 144'h045ff6d9f0fcf5a208bdf7a700230426f82c;
mem[1082] = 144'hff83ff35ff5a042804500a81fc7a052cf16b;
mem[1083] = 144'h0854f0e3f63c0bb20990f7410a0afdb2fb4b;
mem[1084] = 144'hf6dc0831ffa507da0395fa52fd74f8560407;
mem[1085] = 144'h0393faff071cf641f3a001e308c90b260f55;
mem[1086] = 144'hf843fce1f40502cafd5004580d4efc1ff31a;
mem[1087] = 144'hf49afb940b64fcbdfdb0f123facaf32af7b4;
mem[1088] = 144'hfa07f96a04d3060b05b501000a60f2b707fa;
mem[1089] = 144'hf83cfa23f333f4080445f61201edf2170ae4;
mem[1090] = 144'hfbb6f1ccf11c08250a45f56bff0304b507c1;
mem[1091] = 144'hf0400177fe77f2a6f828011a09f1f2300c70;
mem[1092] = 144'h013702c9f5860206f22304b2fd08fce0f65d;
mem[1093] = 144'hf26ef394f9750c6ff8de0319ff3c0880f177;
mem[1094] = 144'h0ae7f4b2f8cf004c06490eebfaeb0ab90c7b;
mem[1095] = 144'h069ff82302abfcf7019bfaa7f5770b51fe29;
mem[1096] = 144'h0e0b0a6df23f0961ff5403f40550ff1601cd;
mem[1097] = 144'h0e02fcab035df86ff27b0797ff1003faf15d;
mem[1098] = 144'hf326fc580f51f8e1f89c071bfe1c087ffd1e;
mem[1099] = 144'hf5f9f9abfa750a8701bdfc3f0166058afc6d;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule