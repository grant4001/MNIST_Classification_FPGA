`timescale 1ns/1ns

module wt_mem0 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h005703bff1b703ebfb39f89aed67ebc906c3;
mem[1] = 144'h02f6f6f600e8f188f28bfc9f073bf367f740;
mem[2] = 144'hf8caf0d7fa98ef75f33def42f4d4f5640901;
mem[3] = 144'hf486fc0dfa35f268f785f1fcf5e40c4b0a51;
mem[4] = 144'h0590f3cefc36ff3408eaf0e5f2feedf40b65;
mem[5] = 144'hed8b0341f93efde9f42b0a220860fa14f213;
mem[6] = 144'h01ca037c037d0bcff642eee8f4f802c4f5a6;
mem[7] = 144'hf8be025afe5bf21cfd29018b0c140272feea;
mem[8] = 144'h05e60d0400b5f324feacf1a7091d0905f346;
mem[9] = 144'hefedf38df781f311eed2ffb8f1a1010a035b;
mem[10] = 144'hf42fffbbf41dfa5ff8d90aceef89f3a0039e;
mem[11] = 144'h096ef07d08510741f0e50c740533f18a0304;
mem[12] = 144'hee47025eef76f602f12fecc9065bf1f1fb8b;
mem[13] = 144'h0bb705880576fb3604a0f0adf3ab040902fa;
mem[14] = 144'hedfd041404e4faa1f9c2ffe4f31d08f7f23b;
mem[15] = 144'hf956ffdcfeeaff70fecbf0c5055700620496;
mem[16] = 144'hf52e0257f8ab08b0ffaa02cff00405ee05b1;
mem[17] = 144'hf4d9edbd06ceefa407a5f82af64aeed9edff;
mem[18] = 144'h0276f0370b6ef44afb24081b024802b4fc26;
mem[19] = 144'hedd1f3f5ec86ef99ea40ee34f4d2fc33ff58;
mem[20] = 144'h013bfeb5006efb22f044eeedf2d50188ee8c;
mem[21] = 144'heeb2f306f1f7f87eeb9af467ec3af231f1cd;
mem[22] = 144'h00d0f65f0643fe73fd58fff2fad4050204b6;
mem[23] = 144'hf5090ab9f3830426ff93ef34f447ff5cf4a3;
mem[24] = 144'hf8c7093a0cdcfdfbf79fefa5043a02230015;
mem[25] = 144'hf3930874f207f3a2fb780b3cf764f9caf9e9;
mem[26] = 144'hf7980bfdee6f06edf18500c80e75f5dff157;
mem[27] = 144'h05ff0835fdd503cbf78cf8d9084ff7f408c3;
mem[28] = 144'heefbf88c03dbf506f60e0d32fb4e0c88fcb3;
mem[29] = 144'h0799f5c90d540da004e30dacf3f0fac90331;
mem[30] = 144'hef88fd1a07d0fb8805e4ed5afa7e02a0f292;
mem[31] = 144'hfee50344f94bfbb40515f89bf26df8b5f333;
mem[32] = 144'h01420247ee79fe7df14b0d63f8d7f33c0c88;
mem[33] = 144'h06a8fc67ff9d0b22f9890024f278f2cef37d;
mem[34] = 144'h08e1fabdf536fe04f7ac0ad409a7fcb9fada;
mem[35] = 144'h0a0107cdfac3f490f4e403eaf5e8ee6ef5e4;
mem[36] = 144'hf597f0cb08cf02980d5808420830ecf2ede7;
mem[37] = 144'h057bee3903bb01acf61bfb5c0c7c0daf031f;
mem[38] = 144'hfc07faf8067803f6fdc0eeacf74f0999f5ca;
mem[39] = 144'h0b57003bfe00f3cffa68030804d3fcca045d;
mem[40] = 144'h0c93fdcf09560ccf0934085cee2ef5b60279;
mem[41] = 144'hf63eee64063af62d03560df506030109f9fd;
mem[42] = 144'hfbf90b37f428f8630064fb0502b9f5a9ee8a;
mem[43] = 144'hf892f23bf41705750af6fc9a0222002408f3;
mem[44] = 144'hfcac000af00cf7f9ff15f770f1d20458f0f4;
mem[45] = 144'hf4f5fa7afb26f9d8f1a7f54706b2faaee98f;
mem[46] = 144'h0791f802f088fdb60dd3066b0908f77e0919;
mem[47] = 144'h0887f08ff9070e0cf8c70ce40a7ef6bdffb1;
mem[48] = 144'h0bb0f59c0891fd36f160065ffe57edd5f2d0;
mem[49] = 144'hf382011ef72b0de0f334f258f113f471fc83;
mem[50] = 144'h0ab00591efa200bbf98efca50414f5740211;
mem[51] = 144'h0b8ff20cf4b4f0d6f643f126fdb70aa8ff5a;
mem[52] = 144'h0184051cf118022c0698f901029dfcfb0614;
mem[53] = 144'hfd0d0474f003f863ff73f7cdf9120085fc5e;
mem[54] = 144'hf49df254ed9ff2e0f3650c02f22c0bfaee8e;
mem[55] = 144'hff130d91fd41fa8d00acfc1afcf70b36068b;
mem[56] = 144'h00d907feef4afb25f334f3e3f64dfeaefdd7;
mem[57] = 144'hf2caf782f4b501480ea503e90d95fa0c0d9f;
mem[58] = 144'hfd6af63dfa52fdb70b6107c00d57ef95fa06;
mem[59] = 144'h0f2d03540a590eec0672f546f764ff72f312;
mem[60] = 144'hf399ead6f261eb6ffdfbff940152f8e1f6b4;
mem[61] = 144'hf29df81ffbe8f10aeb54f641ed59fe670367;
mem[62] = 144'h091ef6ee0983fc67fe93031c075efa4a082b;
mem[63] = 144'h06aeeef7ee43fecd01bef12ef56aef0ffc10;
mem[64] = 144'hed9ffcb90021fa680948ed13f5bbf5c2f0d0;
mem[65] = 144'hfbd801270076010b0577f565f87bfec30742;
mem[66] = 144'hf4cbf715f1b2fb7dfa17051a0c20fdf40d46;
mem[67] = 144'h0be40186fbfffeb00005f2880231f82afdaa;
mem[68] = 144'h0664072bf5fdf922f5940daaf9aefee9050e;
mem[69] = 144'h01b40e6a0ee3ffb40475096bf0cd09450962;
mem[70] = 144'h00a10501fc1df3f4f18ff2f4f74008c6ff2e;
mem[71] = 144'hf240f05b0c67040cf70a0fe20768f74bf8a0;
mem[72] = 144'h01160ed7fd5dfe080f30fb5bfbc403a00b6d;
mem[73] = 144'h0f70027ff35df781f78b0ceaf956fc090306;
mem[74] = 144'h08c2f6c806b8fe2c0af9f00bf440f2210cba;
mem[75] = 144'hf18c0e23061b0ebbfc0a0efd0ae308fdf728;
mem[76] = 144'hfc3df8340b2ef534fe40099d0192fb61054c;
mem[77] = 144'hf6a0f0a0faf2f76c0dafffb3fe1eefdb0d67;
mem[78] = 144'hf556f5620312fd4f0bebf6e5f7940fb5ff75;
mem[79] = 144'h00e107b4f4e707d305c4f52b0e480458f4b5;
mem[80] = 144'h0d65fd3907c6fdbd0fb10943f8d10dfa05ec;
mem[81] = 144'hf92c03840c6df022f4adfd24fc75fa49f5d8;
mem[82] = 144'h064af2acf852f3ff0fce032e01d9fa4403ae;
mem[83] = 144'hf4910c1a009208e007920787f631f1bb04f4;
mem[84] = 144'hfb41fd03f57a03ed0e6bf30808a50a9cf5aa;
mem[85] = 144'h0f760eb3f8fffacc0cf20f1105810e65f0c4;
mem[86] = 144'h08b700aef20d0582f904f67206a6fb2b06ab;
mem[87] = 144'hf082f9fc0d5a01670d680383f0f0f47c0d34;
mem[88] = 144'hfcb8fd29f3c3fac3f0edf3e1f09d01630b0d;
mem[89] = 144'h0104fb17f7e2f65c036af5410b91f69ffffd;
mem[90] = 144'h0462ffcd07500031fe9b0007027dfc39f2fc;
mem[91] = 144'hfc71fa7806c805c40b090a00f04dfe770ef3;
mem[92] = 144'hf80ff14cf6acf625f8810c0f068d0033f31a;
mem[93] = 144'h0fa5f66804a7087700a1fcedff41f9900511;
mem[94] = 144'hf6b90bd40e370925f23cf38a0b270d820ed0;
mem[95] = 144'h0fd6f8ccfd94f09bf87af6c0f1620c730b08;
mem[96] = 144'hf618f3d0f7ebf8bffcda0747fa160510fe82;
mem[97] = 144'h02d00f630f3e078df03bf65a07abf8aefd61;
mem[98] = 144'hf420f25402d803a60f79f7430813f42df2bf;
mem[99] = 144'hf66b0f9ff2ee09fbf3960a53068904e602d2;
mem[100] = 144'hffa7f5f6059bf5d00f47fd49003b0cbb03ec;
mem[101] = 144'h0119f741f28f080a09c107bb05a807bb0feb;
mem[102] = 144'hfc61f8240d090d3ff449f0cafb3e06a40621;
mem[103] = 144'hffca0bbb046c03170c77f085f34806c6fef1;
mem[104] = 144'h03150bb2f8b7fa59f3fef8380dca0d8f0a23;
mem[105] = 144'h043904840c50005a0a55faf60cc5f5b4fd35;
mem[106] = 144'hf18806e7f733faed09a30bf80358fcd7f2d8;
mem[107] = 144'h03760fb705adfced079a03fb0c6b08f7f2be;
mem[108] = 144'hff350d480548fdbffa9bfa210e59f2f3f519;
mem[109] = 144'hfe10f92402caff7d049a0d9a0a35f14e0266;
mem[110] = 144'hfca001fffd4bff8108810336f8f7fc9d077c;
mem[111] = 144'h07c90d6fffdb04cf019300540851f9200d9a;
mem[112] = 144'h094e05250b1df72c0ffa04ea0cf200540ae2;
mem[113] = 144'hfff30eac0a610ccbf464f80a0c87f21afe62;
mem[114] = 144'h0e450865ff1efb330edd06d60c98f4430416;
mem[115] = 144'h03def0640ce7040b0c43fafc04d7f8de07d7;
mem[116] = 144'hf916f1a5fccb0dabf810fa54039a00390bf1;
mem[117] = 144'h0485f844f4a106830342f8e8fbfcf1bff8e9;
mem[118] = 144'hf13c055c0f05fac6fe9005c90698fa920723;
mem[119] = 144'hf6bff554fc7009be0c7f0cde0c08f8de0f54;
mem[120] = 144'hfade0d40f197f31cf100fc92f6e1f6a50290;
mem[121] = 144'hfb36092f0619046505eaff26f2400745ff87;
mem[122] = 144'hf956fdc205db0f52fc12f91e0917ff49031f;
mem[123] = 144'h0ba50ef40477f3e301d8f30705610957f9c9;
mem[124] = 144'hfa56fadb0d2ffd09f6fb0648fcd001dffdfb;
mem[125] = 144'hf6b0f605fce1f1bc0e7508fefe56fb0f0a99;
mem[126] = 144'heff6f6b9fa730bdffec7f5f60552fd9ff76c;
mem[127] = 144'h0bc6080bf06df77102d2feab058e00a70b62;
mem[128] = 144'hf8d401c7ff6f00b50bfb0f3f0a490d340224;
mem[129] = 144'hfbf7fa16fde9052af1fd0967fb4803450f2b;
mem[130] = 144'h0c5d0a29f65bfb9c0552072f0ac409a5f5fc;
mem[131] = 144'h08ccfb26f684fb9600e8f457fa92068b0454;
mem[132] = 144'hf8820e330ddb06d8f91b0b1405f80aabf5b3;
mem[133] = 144'hfac5fc47f532fdf90b5b06dafdcdf60b088d;
mem[134] = 144'h0f730b5f064af698f733078902af038efe17;
mem[135] = 144'h09a80ba20e2500aff8fb0924fa7f0227f2ca;
mem[136] = 144'hf6190929f0a80058f7080f38f2c20a7b0f8d;
mem[137] = 144'h0f73f6daf7aaf42af158fb270bb408460d73;
mem[138] = 144'h017c0cfc0845059e01dbf8b20b78f6c00899;
mem[139] = 144'h01c308350c2ffec6f81b09570c1bf8d8f5bc;
mem[140] = 144'hf9b80412fbd6f997f7500d8b0be50267013c;
mem[141] = 144'h0d530147f85cf5580a4104fbf75ef5daf26f;
mem[142] = 144'h02c50ac90813f7f60e920aa90af4f3ad04bb;
mem[143] = 144'h095909bbf9040f290e81f0710cc8f2c70332;
mem[144] = 144'h0bd9fdb10edefbf204a7f80b0aedfab2f7b5;
mem[145] = 144'h0f3e0f560938f43c0833fd21f8150b820baf;
mem[146] = 144'h007a07b1f7a5f231073cfb03f42f00ca08dc;
mem[147] = 144'hf7e5011bfc390c66f02d054e00b0f427001b;
mem[148] = 144'h087afd75ff3d0aa20ad30e55f2af022a04a8;
mem[149] = 144'h0f6f0c05013b0a4af504f323010d07e2f103;
mem[150] = 144'h00bbff1ef7de025b01a0f4c7f368fea7fa7e;
mem[151] = 144'h023605240395f33bfa0200450f68f33f0351;
mem[152] = 144'hf029fb0a037df16cf45efaa3017afc48f804;
mem[153] = 144'hf4290eda0bfaf86805e202730d830f4000d8;
mem[154] = 144'h0ceafe7ffb33f60efce3ff3f01310a290b5f;
mem[155] = 144'hf7e2f4fff1900e6df49008aa01e20ba2029a;
mem[156] = 144'hf5f10ed2f16bf306fc110c77f214004409cd;
mem[157] = 144'hf37bfefef4610fc6f8cb0ca5ff26f8dcf56c;
mem[158] = 144'hf5280d8c01a4f707ff04fdcc02af0d7bf51b;
mem[159] = 144'h0770faa9060d0c1f0b84046a08070b3f0198;
mem[160] = 144'hf40afeeafc92f3160293fe98fdd1028cf239;
mem[161] = 144'hf472f82dfcd207dc053c0bfe03d1f9700a81;
mem[162] = 144'h05bd083b08d70bb7fab0f10cf60d0e320ba9;
mem[163] = 144'hfbd107dc04f5f7daf5140a85f0ca00bd0df8;
mem[164] = 144'h02b3030dfcdfffe309aa075506d008c20c4a;
mem[165] = 144'h0c5a0eb0fef30a02fa290d1ff1a8f36e0b9e;
mem[166] = 144'h0af10cfb05620120f20df9cd048bf6d10146;
mem[167] = 144'hfa5ff3590b1105b5007b080202cc0e18f10c;
mem[168] = 144'hf433f21a0dd50066084301befdb1087607c4;
mem[169] = 144'hf89bf5e6072406d80c9101be0c9905ae08f3;
mem[170] = 144'h0699fd8df7a5f7a80789f31803360dd80a51;
mem[171] = 144'h042309f3f0d00c63f197fcc707fd0fc60251;
mem[172] = 144'hff76f042feacf76208e9032c0988fd58f833;
mem[173] = 144'hffabfafc06ab092df49604880b67f457f5f8;
mem[174] = 144'h0039f904f8cb00c0f1570735f1f00382f0ae;
mem[175] = 144'hf9f3f2350d79038cfdfbf4a9f772082d0019;
mem[176] = 144'hf9410b93f6fefe3af3fdf24cf87dfb3a0cb0;
mem[177] = 144'hfff6fe40090809acf2abf2d10c9a0f7804be;
mem[178] = 144'h0f410e870391fea700b60afdf4c10f64fa70;
mem[179] = 144'hfae10ecf0809f1f4f8540582f099f13b0322;
mem[180] = 144'h012f0067f6140ed2fbd605e2f97af9fef804;
mem[181] = 144'hf36a041cf8410a0b0031090ef7310f05078b;
mem[182] = 144'h0c4ff1c3f2a4fbeef314fa940729fd940b25;
mem[183] = 144'h006c0f1bf5930a0b0d69036bf83afb87f92d;
mem[184] = 144'h00fd083306f2f12af17e088b00b3f6b2f9b3;
mem[185] = 144'h074d05fb06fcffe1f1d70ead05530a19f2c3;
mem[186] = 144'h0f6effaef6e9f2fb093605c8f4140ba2f931;
mem[187] = 144'h00020f2af05ef8b3f960f503f6170979f86b;
mem[188] = 144'hffb0fcfe067a07520084f3b7fa90feb400a6;
mem[189] = 144'hf19ff657fe4fffc30aa3fd10040af81dffa7;
mem[190] = 144'h00f2ffb50282f235f38ef5ff0005fa280b8e;
mem[191] = 144'h050bfa17fe20f2850883f1b10bfd0acaf075;
mem[192] = 144'h06b80e5a049a0d440d970d7008860668f3e7;
mem[193] = 144'h05480de80c62095ffac5f308fe1efc780d1e;
mem[194] = 144'hf403fedef496f278f8bf08a6f0eafd17f452;
mem[195] = 144'hfe96062df5720730f136f475098cf3370463;
mem[196] = 144'h0faf0ca9fac90afcfb9c0486f774f37102c2;
mem[197] = 144'h03d9f8ea058dfffbfc7ff4d9fd9908a2f368;
mem[198] = 144'h05daff700eccf293fa45f5f60b8c04490d0e;
mem[199] = 144'hfd2ef6880d34fc080113fd6ffb2b042bff5d;
mem[200] = 144'hf4f702f3f170fc25f6ae019a0c8b0c1bf07d;
mem[201] = 144'hfea60c0504f0f511f2feff68fc05f500f31c;
mem[202] = 144'hfc8eff06f7ca048404dc0c41f4a2ff3f05d9;
mem[203] = 144'hf442fcbbfd5cf99bfca2f7a70e7cf4a4f412;
mem[204] = 144'hf9560c5f0dc3071ff474f46d08c1f53ef73d;
mem[205] = 144'hfb66fbee0af00799023ff8e90c90fb7af992;
mem[206] = 144'h0897fd8d0c18fd26f6b1f63e0038019ef4fa;
mem[207] = 144'hf076eff6080609170184f01ff51fff3af771;
mem[208] = 144'h085cf2a6fe62fb3af9f90fe3041906ff0155;
mem[209] = 144'h0b43fa9cfa7b08c6fad2f82c04200b1bf033;
mem[210] = 144'h0812092d06ca0cda06df0040f049fbd20861;
mem[211] = 144'hf577f8b90081087905b7fc04f372feee065b;
mem[212] = 144'h089af5e3fe16f3a0f8aefa1afa1c0623ff91;
mem[213] = 144'h0be0f2f9f3cdf50bf8eefd47f4910fd00b8d;
mem[214] = 144'h008f0d3c0531fd4403ee05d2f09d0a7603d4;
mem[215] = 144'h013e0138f508efd90592f7d1ff810ee0f563;
mem[216] = 144'hfda101f00b6002800f1af91bf233fe3af8b8;
mem[217] = 144'h0af00ea20664fb65fcb1ff0bf6f8f24ff87b;
mem[218] = 144'h01ff04c007530f130f690d5cff080f14f3f0;
mem[219] = 144'hf6c8f3730904f612022afbe4f0a901b70567;
mem[220] = 144'h09e10be7f6d6f356040bfb22f1d9fef50a7b;
mem[221] = 144'hf73af1c1f115f478fd3df03d07a40073fc0c;
mem[222] = 144'hfc6e00befaa309f30930f7c4f4a8f7490904;
mem[223] = 144'hfb580c4e02540e2df6c6f0410a8c07e5f2d0;
mem[224] = 144'h06ad00e7f5aa026e0dc3fca1f6b807cdf134;
mem[225] = 144'h0e2f0085f03ef5a8fff8f1500050fa6bf8e5;
mem[226] = 144'h0a77fd85fcd9f90308e5069f0316f742fa32;
mem[227] = 144'h07dc0e6f0fd90cbff0e605b5060a06bd0b8c;
mem[228] = 144'h02c1f2fdf46a0df5f84d076df90607bc0ad9;
mem[229] = 144'h02d7f679f80e02b00c6e0e8e0f9efa270a49;
mem[230] = 144'hfe24ffacf39f0485080e0211f4d606ad008c;
mem[231] = 144'h0f05f09cf433f085f399f69af8da0119037c;
mem[232] = 144'h0d7d05e4f19c0df1f89aff72f2770c9d0fb9;
mem[233] = 144'h0f97fe56f024f3dc0c9e01e2fbfbff490e51;
mem[234] = 144'hf945ff2809bd05990f730ed40738f5ee04df;
mem[235] = 144'hf61a019f0e6bfc940f81faf4f2c0f941f76e;
mem[236] = 144'h073009eff7c5fce6087ef2550269fcc70b97;
mem[237] = 144'h0919f008f999f1500be9f6c1fbf3fc5903ce;
mem[238] = 144'hf37c0f4cf8da0dd7f787f06307e3f525f2b6;
mem[239] = 144'h0210fb81f3e6f25c0362f8a3f050f9b209aa;
mem[240] = 144'h0632f264f510f403fe1df0c8fec20357028a;
mem[241] = 144'h0ac20390f4ccfe2ef298f255f8ff0ef9f018;
mem[242] = 144'h09010e33fecb03a4f2980951037dfe43f812;
mem[243] = 144'hf3220d0b0692086bfff1008208cd033dfc26;
mem[244] = 144'h094ef1cf0f5e06070fd2f50bf804fcb3f1a7;
mem[245] = 144'h087f07cb02da0d17f9bbf6090b23077ceff3;
mem[246] = 144'hfc2aff64f274f3d2fe0f014f00cbf59200fa;
mem[247] = 144'hf248026bf8ccf84c0367fa540994f1070021;
mem[248] = 144'h0a7604080a02f088fc5a054bf64bfb50fbf3;
mem[249] = 144'h0be1051d0ab906f10557064002a0fba50f00;
mem[250] = 144'hf7adfffe08b40154fe300ba207c90363f8b9;
mem[251] = 144'h01e50466fe460edff8bff7e602040bf1f116;
mem[252] = 144'hf576feabf86a0f1bfe7effd301970fcf0269;
mem[253] = 144'hfc71f6aaf286f4caf07bfe9504a1fd8bf452;
mem[254] = 144'h063e0c8ef2000e4a0d4bfe070d78f220f776;
mem[255] = 144'h063af4c00816f3baf3c806f3f0e4f84cf725;
mem[256] = 144'h0cca0a1503cef3fc05d50bec07dff4a804ec;
mem[257] = 144'h0084fad807070a03015afb0801b103a0f473;
mem[258] = 144'hf61befff06970525f70cfa940d65f860f65e;
mem[259] = 144'h0c7dfe89f2790e30ff450f3b094af66f069b;
mem[260] = 144'h0190f184fe11f9d2f17a0852f3e8fb1707a9;
mem[261] = 144'h07ed05d0fb2bf93e0a54f8a10db20a0404ed;
mem[262] = 144'hf0edf897f0f605acf7340dbdf70a0253f4ea;
mem[263] = 144'hf150fdbffae80dfbf8c3fb3bf859fa9e090f;
mem[264] = 144'h0f7c07a4f9c5f9f0f1d90e59044f060c0f90;
mem[265] = 144'hfcbff59603b4f88e0a330c96f7c304b906e2;
mem[266] = 144'h06e50395f50a02c70f380caafb05fe700e6a;
mem[267] = 144'h082b0946f30c025a0fdef88bf0c2083ef120;
mem[268] = 144'hf9c5f74ef5ad0c810476f219095ff6ba0ead;
mem[269] = 144'hf56f0582f65d08080a590971f21afb76f8c0;
mem[270] = 144'hff0c0e7f059300c2fc690172f4aa0deef57e;
mem[271] = 144'hff1efc97fc4006390379087bfbb3f7b70875;
mem[272] = 144'h069bf041fdcfff660766fa1e0825fb00f5a8;
mem[273] = 144'h0e7b02dbff7afb8efa58074402a10d77014d;
mem[274] = 144'hfdb00f2ffc9af62af64b0d2d0777feaef231;
mem[275] = 144'hf299075bf13c0108f8bcf87906b303ca00b9;
mem[276] = 144'hf26e05b1097d0b7a05a1f2f0055df18201b8;
mem[277] = 144'hf40a00ed008afb19f59ff17e0bcbfd1d0407;
mem[278] = 144'hf6c4f2b5020c0a5101e2f0c90ae608baf425;
mem[279] = 144'hf896f5eff2bdfcccf39afcd7f5dbf273f447;
mem[280] = 144'h0b3d07030bd304daf65a0cd6fa270299f823;
mem[281] = 144'hf9ac020bf937057f0b8ef8cc0db208d60525;
mem[282] = 144'h007b0767faf606640afaff9af1dbf63dfd30;
mem[283] = 144'h04faf1a70dfcf02e02d6f703029407e80e8d;
mem[284] = 144'h05db0488fc890fac0b7b0723fc15fa21fc80;
mem[285] = 144'h074efda2f37af873f662f35e09f9fd03f8f5;
mem[286] = 144'h0de5f708f32befdd008cfd4bfb3103ec0b4c;
mem[287] = 144'h083ef4840e7cf4e7f113f04d03f3f42904ab;
mem[288] = 144'h090df87c043608cd0b420b6601bdf0b1ffd2;
mem[289] = 144'h041af6f600fb09baf37601bc0d7efb84f58f;
mem[290] = 144'hf076023ef05b0eb603f80274f9a2fdda01a9;
mem[291] = 144'h090201d7ff9b0e9d02d20bb50e4a065ffba1;
mem[292] = 144'hff2dff2b0a2a0e59000d0ef7f8e3fbf9fdbe;
mem[293] = 144'h04600accfab7fa730b2af4b1fca0fe4af694;
mem[294] = 144'hf2b9052d0ab30b3bf6b80526fdb4082802e0;
mem[295] = 144'h03b70dc6f625f4cc0bf1007107c40933faf8;
mem[296] = 144'hf668faa8009bfa940af50b1af33b0a0d04af;
mem[297] = 144'h02ce0c0201d9058c041f0671fd6803ef0b8b;
mem[298] = 144'hf0d1ff21f0daf39ef110f763fd55f9b5029e;
mem[299] = 144'h06bafbbf0c440d5aff6bf0db0be40e43fc88;
mem[300] = 144'hfb49f5d2f2f2fcbcf56007c70101f8e70c21;
mem[301] = 144'hf1260f53f66ff4f1f4ab05aaf1ee09b4fd95;
mem[302] = 144'hf4d7f3f00ac6fb00fc55054bf91bfbe0fc44;
mem[303] = 144'h0735f1e3f1a00ebb0729fec3ffcbfdb0fbc9;
mem[304] = 144'hfaa006b90281ff9df72a0b3d0a80fa49f02a;
mem[305] = 144'hf82efb250bef09ecf4080535fb42f089f217;
mem[306] = 144'hfa68fb14f25705480733f936ffb4f813fcc4;
mem[307] = 144'h0b270fa6fe200f1ff904fbe1f96af9d9fdb5;
mem[308] = 144'h0b300da8f76805d1f3a0037cf7dffbbd08f3;
mem[309] = 144'h0ceafeebf0b70744f97af26cfc080254fdc6;
mem[310] = 144'h0963f3de0882032df89e08bbf95af7d60352;
mem[311] = 144'hfcb009d7fa67f9bb05640d1405befce4f4a3;
mem[312] = 144'hfa6df82fff4ffae003c0086901bcf52306e7;
mem[313] = 144'h09a6f60bf389f85b025203d904cff148fdaf;
mem[314] = 144'h0cf2091ff0eff2eafd5dfbebfef0f9f10651;
mem[315] = 144'h01720c4cfebef8260f25f2ee0cc3022201e8;
mem[316] = 144'hf442f6b1f48ff36b03c2fd8d0e2ef874f12b;
mem[317] = 144'h00950fc50e0af8b4fd20f55a09e3f49c0d25;
mem[318] = 144'hf0950565023ef59c06e8f8f401ba08aa0268;
mem[319] = 144'hfb7cf0070be20544fa9f0904f2690cc20cd6;
mem[320] = 144'hf6160c39f123044a0d90060df5e900f70571;
mem[321] = 144'h092309aaf2870b96fce2f5dbfb0600600975;
mem[322] = 144'hf44c01b302b301170a78f869f840f43a07ce;
mem[323] = 144'hfe69fc69ff8600aa0d65f4550fdb09ba05eb;
mem[324] = 144'hfce3fd19046601edfeba0ca3022df8e9fca0;
mem[325] = 144'hfaaefa48fc9f061cf0c30692f0ce084c0da8;
mem[326] = 144'hfcc2f3520fca097cf571049c0269facd0461;
mem[327] = 144'h0662051f0873f511f460f3810631f3efff65;
mem[328] = 144'h0addf747fe3908e8073af420fd97f52106be;
mem[329] = 144'h033f006df6e1ff37fe6bf8f0f139017df81a;
mem[330] = 144'hf70300a2ff4403f70ea3f5e0f1cf0354f92c;
mem[331] = 144'h01b105e1ff55fe3e0e41f28702f6f31aefd7;
mem[332] = 144'hf4fff43a0be90dea0214fe33f3c7051bf981;
mem[333] = 144'hfbd4f24ef862f3260accff030e9606490296;
mem[334] = 144'h096a0a62059effd40d5a0c3ffcccf1ee058e;
mem[335] = 144'hf9b402c80a5efd900874fa8b085afc7c09de;
mem[336] = 144'hff2b07b8080af9670efd0ce3ff08f1a501c7;
mem[337] = 144'hf2c4fc4deffdf5c2faabfb10f37d0c49047a;
mem[338] = 144'hfe6af995fe300bc9f09a0c7c0773fd68ff96;
mem[339] = 144'h035e0c31f5390afaf02cf2a501bef5b0f73d;
mem[340] = 144'hf7930bd5f83ef4cc06fff636f1a40d41fb6d;
mem[341] = 144'hffb502ca0024f8cdfbd8f23d08ca03c6fe9c;
mem[342] = 144'hf194fe130339071208c70f82fb030752f1df;
mem[343] = 144'hfc57f99c0d05fbf908ecf5b3f530069bfeef;
mem[344] = 144'hf2200dc3facef741f477052106aa01f2076c;
mem[345] = 144'h0ba6fd330122ff52fe130d02fb0c0a42fd96;
mem[346] = 144'hf8940fb4f0aa0c4909e0faab0417fee2f449;
mem[347] = 144'hfa67022f0531fae1fe190e070cfd02f5f03f;
mem[348] = 144'h066d0fcffb02fc24f522031dfb88f83afbae;
mem[349] = 144'h080effc9f4d2f3560a39f1bb02b3089f03ae;
mem[350] = 144'hf340f690000204ee05480a070d470dddfa95;
mem[351] = 144'h063af3c50b12064b0e2408a1fe8f0b870013;
mem[352] = 144'h09bcffd202390f4af6650bf00f2afe500f0c;
mem[353] = 144'h058f04800471020af987f4740868f2f20d8b;
mem[354] = 144'h0250f50f0da301d3f677fbb7f3bc0032fc50;
mem[355] = 144'hfb570c85fb6c0ca201ff07a404fef7b80f52;
mem[356] = 144'h015306b8f3f80f8f0ebd0f9e0a57051f051a;
mem[357] = 144'hf7360477f4250bbffc5300b1fb45fa09f371;
mem[358] = 144'hfa0f0195fbb6066df2920e770b5bf91af1f5;
mem[359] = 144'hf404f1d2fb400541fc73ff02fc54052b0ae4;
mem[360] = 144'h0981fe48fca1f2020f8c030e04ec0241f381;
mem[361] = 144'h0e4ffc81032efd02f2bd091df96a00c40b41;
mem[362] = 144'h09c604be0beaf442f96200b2fc1bfbdc0b90;
mem[363] = 144'h0eec0e0f0d2ffc8bfaa40333079f0de3f72e;
mem[364] = 144'h0eca0a100c1af637092bf957f47d0327f334;
mem[365] = 144'hf8b50f6404fb00a60fb80469f6420da80316;
mem[366] = 144'hffe90588f1f7f035ff7507aafd270cbb0d70;
mem[367] = 144'hfd21f0b9f94a0e540841fd63f6a50aa5f86c;
mem[368] = 144'hfa08f62df1d10f1ff5d40ae200d2f4dcf373;
mem[369] = 144'h0324fc910aefffcb0bc908fa04f700c0f83f;
mem[370] = 144'h09580549f305f0aefedaf4cc07dffa60f1f7;
mem[371] = 144'h084afc5a0c2e0dccfbc7fbe30e4003080f37;
mem[372] = 144'hfbce0e27fd060a1400ecf7b8f12efd9dfc9d;
mem[373] = 144'h0872f08f039cf2ba0b6808c5f65609a605b6;
mem[374] = 144'h0be10ecdf08a0e04018207d8f92bfe340352;
mem[375] = 144'hfb64f23efc6c0769fa13f9fd0455f8eb010b;
mem[376] = 144'h06c20846fc770df7057ffdce0e640bfcf454;
mem[377] = 144'hfa5cfebf0c5c0bcff0ef0df4f9dc0f2f099b;
mem[378] = 144'hf20a012205b504f4f7310935fa930e09f9d6;
mem[379] = 144'hf3a1f9cc003df996ffe5054f060a0ed50f86;
mem[380] = 144'h0b2a04f6fa90fe8bfc50053f02d50650f48b;
mem[381] = 144'hf34a0243fd4bf6a0056bf7a601b30d76f07a;
mem[382] = 144'hf12a0ae70b240432093e0849faa7ff32078f;
mem[383] = 144'h0e5702b30c7ff745ff310beefec30258004e;
mem[384] = 144'hfa45fa0af739f51d0b8609a9fa9906faf1cf;
mem[385] = 144'hf5b8f49f056f03eb0e7100f7f68902c9f3fe;
mem[386] = 144'hfd6e05dafbe3ff72fbfb0e4109e905e8f6d6;
mem[387] = 144'h02dc073c07bffe83fbb1fc01f7300bc8f943;
mem[388] = 144'h0845ff5cf22a0d300deef726f88c0400f5b6;
mem[389] = 144'hfcf4f12c0ed4f22f0d81f215060e08690ef2;
mem[390] = 144'h0dca0231f77df5f90742f2e1fe1c0ae4fd1b;
mem[391] = 144'h0ad10580f514f4510b8e0dd2f4e5ffca0a27;
mem[392] = 144'hfb6bfd2a02f3f1e00c8c071b01bb031102bf;
mem[393] = 144'h0ef00af1f4d10bfe09d40c84f36701030c80;
mem[394] = 144'hf63e08ba0a1b09dcf581031b03fe0d320ae4;
mem[395] = 144'h056f099207edf101026b088e082b04f6fb7e;
mem[396] = 144'hfb5e02bd0a15f38c0b3cf3820175fdb7f47b;
mem[397] = 144'hfc05fb40035ff3a3f2e0f6cefac70502f765;
mem[398] = 144'hffe70eba00edf929f027fe0706c9f2cbfba6;
mem[399] = 144'hf263fe580167f190055e099b0e6e024afac1;
mem[400] = 144'hf4acfa96f01ef32d08b901cef836067903f9;
mem[401] = 144'h011ffc6cf67c09ebff3dfd260050fcc1f396;
mem[402] = 144'h010a0953017309d3fade04d307a1fdf2012c;
mem[403] = 144'h03880d10fd3c0828f099f9a60f4909f6fa98;
mem[404] = 144'h0897fde1f37705df0faafcddf990030ff1ba;
mem[405] = 144'h0eb9f1c0f2af0edcf80b050df6aaf7a6fdbd;
mem[406] = 144'hfd6bf24305970cc404c5fefd084a0f38fdcc;
mem[407] = 144'h06e701510af2f7c00d170becf52707b2081c;
mem[408] = 144'hfd050691f2ddf1b5f7ac0e88f2d0ffe6005f;
mem[409] = 144'h008ef33f0fa7fb8d0579fa990b630e03f42a;
mem[410] = 144'hfda7fcbbf6250170fc50f217fa650eb40122;
mem[411] = 144'h0c23fc68f602012a0ec4058209200b2af2cb;
mem[412] = 144'h032202df0d64faed0c33f375fa84f0d30d7b;
mem[413] = 144'h067dfb37f462086bf51500fef4af05ccf055;
mem[414] = 144'h0b3908a5f8f4f14d0cd902dbfa7c0701f526;
mem[415] = 144'hf6080d400bfbf0f0079b03f70c91fb45f2f8;
mem[416] = 144'h053cf592037cf98c026508120eb40484f0c6;
mem[417] = 144'h07ce0f4e051907ae0153f5cc019502f2f145;
mem[418] = 144'h0d9ffb27f392078df20b0f6efac9fdf0fd24;
mem[419] = 144'h0afb0cee0d090e0a05fdf96cf57502e10fe2;
mem[420] = 144'hfb14006200f2f9b2fee708fd05310f60f7e8;
mem[421] = 144'h0398f20cf9e004000281fdeaf391003df79d;
mem[422] = 144'h0bb7fb99fdba0d8c04e5f355fc4103aaf28a;
mem[423] = 144'h0221ff85f6d10f3ef8b60fa909f6ff03f13f;
mem[424] = 144'hf21c0559fc9100b403b8f1f9fdbcf9b80453;
mem[425] = 144'h077402aef73202b6f8eb03cff0d808ad08c6;
mem[426] = 144'hf0d4f0e5fe9ffd3cf7da05ad0ccc0267f519;
mem[427] = 144'h079b0e3e07930d4e0ef5027f09fe00e90504;
mem[428] = 144'h0b9ffdcaf1650bfc01aef7b8f96d0077083a;
mem[429] = 144'h02fafde509890c5a0c6bf1cef5aff6a8f2dc;
mem[430] = 144'hf2b8f3f306cff824f4a1f20d0154f1fb00c2;
mem[431] = 144'h03d1faeafbf8fca5fb2003d6fd810c1df06e;
mem[432] = 144'h04390fc7066d06da0b490d4b0678f12b013b;
mem[433] = 144'hf6ec0dbef8defd6df6400d69f33ef94a0500;
mem[434] = 144'h0cc5f7e50cca0244085cf63302b209500cc2;
mem[435] = 144'hfe9ff281f2d109c501a8f84c0e1df00e0934;
mem[436] = 144'h0ef300bef6be076afba40ada040308730cda;
mem[437] = 144'hfb50f24800ee0877fa5dfc930e25f4810c2b;
mem[438] = 144'hff4ff065f51606fd05e9fbdff799f574fccd;
mem[439] = 144'hf8cf01f4eff806830b36f6150a300c39f322;
mem[440] = 144'h0ab30d240c8d0f28fd7df8b0f9d2fb600d05;
mem[441] = 144'h048cfd4a0e880996f60afebff4070f6bf993;
mem[442] = 144'h04800b56fe21f8b6ffd4f1ae0944fdadfc89;
mem[443] = 144'h0df1f8260109f8fc0f62ffb204d4f45109fd;
mem[444] = 144'h0a2800a806f9f68e065bfbd2022bf6150ab3;
mem[445] = 144'h0ce9fc9308a6f424f296fef50da2fd0e05fa;
mem[446] = 144'hfb4a026bf28800560819f975f718f3c5f681;
mem[447] = 144'hf6a6f087074201250c89ff5af54afa56f1c9;
mem[448] = 144'hfb860441fd820d1a0854fcf205140bdb00ce;
mem[449] = 144'h02dc0623f67efd21018405ff0f48ff10f7f1;
mem[450] = 144'h016ffb0a042bf014fce00a85ff010a19f1cb;
mem[451] = 144'h0c3ff111f5bf0daa086afecf0e9f0e38096e;
mem[452] = 144'hfb62ff01f0cef8d6f2e4fd1a06cb06fc0f6e;
mem[453] = 144'hf6ab0edffe51f46bfef403460b5df4250e5f;
mem[454] = 144'h0d11fec80122fbbcf34ff223fc9af1eaf361;
mem[455] = 144'h028309a90e9afda9f1f40a010bdcfb49f90c;
mem[456] = 144'hf9770786ffc8f156fc33021a07500a48fb3b;
mem[457] = 144'h05baf8f2f53e07adfc5ef3a909670120f632;
mem[458] = 144'hf0d00be8f7350572fcf8f832f0c9f02cf247;
mem[459] = 144'hfec00219f4160cf4fdcdf88b018e0826f493;
mem[460] = 144'h0b6afa710f53f12f0feff35409ad03de066e;
mem[461] = 144'hf2c80807f51307bef33cf1490860f34701af;
mem[462] = 144'hfd5cfa7cf7cefeaeefeafaca05d5f4c2fe14;
mem[463] = 144'h01e9f93a0110f8daf0cdfc74f572fc5e091d;
mem[464] = 144'hfd39063f0f310ed7f31bf2e2fda1fea3feb8;
mem[465] = 144'h044100de00a40279f52f09f506aef37001a6;
mem[466] = 144'h0cd6fa7c0cd406d50593ffccf2ca0810fe1b;
mem[467] = 144'hffcb02450e32fe2209250f7bf599095a0431;
mem[468] = 144'hf62e0ea10fcb03b00b03fce0f8cb0c18ff7d;
mem[469] = 144'hf274f2a90e0dfa0807a40fb80b9b0521fc5d;
mem[470] = 144'hf7fa0e8002b5064cfb410cfff63505d00fbe;
mem[471] = 144'hfc5c09630f31f498044b039ff3bc08410162;
mem[472] = 144'h0cabfa1c0d17fe730cbe08a8f63d009dfd9e;
mem[473] = 144'hfbc40b440536f66804200dd4fd4e0636fd52;
mem[474] = 144'h023d0db9f36f034009440f7e0b1ef0c6f482;
mem[475] = 144'hf8d90bf000e603100a6704c0005a06560c6e;
mem[476] = 144'hff49f79afa57fc6ff922f5a2fc9af9b306ca;
mem[477] = 144'hfec4f8d3f7affe50fe9b0c1d0823090501ef;
mem[478] = 144'hf0260ba3f4f109eff511f468f334fe41050e;
mem[479] = 144'h0ecdfb8308010bbb058dffd4016d039ef004;
mem[480] = 144'hfb56f35c09cefee8f29f0df40c2a08dd0095;
mem[481] = 144'hfd4f0605f419fed30eb2fca4f432f3eff82a;
mem[482] = 144'hf1a60d85040ffe25018802e50a8309400134;
mem[483] = 144'h03edf049f3360aa5f7d3fc36f1bcfcc609f6;
mem[484] = 144'hf2e50b5e079ff968fd3d08b10fddf054f466;
mem[485] = 144'h02bafe8b06dbefcb053bf3f0f402f23c0857;
mem[486] = 144'h00d80f4109dbf59f02f302f8fe19f7580690;
mem[487] = 144'hf570f3830959fea70c1df76d0454f222f3a7;
mem[488] = 144'hf9af0c31f4e6091d0acff747f50401fa0947;
mem[489] = 144'h0683fa1afa7df5acf6ff00c60e6ffeecf18c;
mem[490] = 144'hfa78034402b00410020009bf027a031703fe;
mem[491] = 144'hff2c05900349f3f7002cfc0200e4f8f70042;
mem[492] = 144'h06290b33fd39f03706b2f8080607f74a0e2f;
mem[493] = 144'hfbf70aaf09d70716f8170e53ffdaff73f00e;
mem[494] = 144'h04370acd0d02fc9af0c2069dfb82f3550eeb;
mem[495] = 144'hfcb708f7f17cfccbf46b0f550bef092df64d;
mem[496] = 144'hf3330120fb5af869fdc302b50405089802d3;
mem[497] = 144'h05e7f211fdb102e0f520f50ef63f08b2028d;
mem[498] = 144'h09e00831f0640502f19ff16b05f3000af440;
mem[499] = 144'h01fdf658fc650f87f6500e19f8950bf3fe53;
mem[500] = 144'hfa06f9c50f6b0094083cf7f8f99d0244005b;
mem[501] = 144'hf8700e99079c01caf1fff646f757f673f332;
mem[502] = 144'hf7d5f493ff070deefb020f3d03c90542fed9;
mem[503] = 144'hf0b7fff9f5d80330f3b7094b01e7f044034a;
mem[504] = 144'hfd00f944f94c0aaf0166ffe1f74507dcf953;
mem[505] = 144'h0188f175006cf7caf1320d2000d2f822f918;
mem[506] = 144'h0f76f66e027bf4a90445f7def2faf438f18c;
mem[507] = 144'h0c4bf7f9fe87f0840293f6b9f006fe63078f;
mem[508] = 144'hf5e40d3d0cc7fa89fc8b0c7f0d14f2c50444;
mem[509] = 144'hfff608e80c3607fff659f13ff509fdea0457;
mem[510] = 144'hfaa4f9e1effdf942fa50f36ff1060a61f055;
mem[511] = 144'h0912f3a3f1c80a7900f5f210f60bfcaff459;
mem[512] = 144'hf9e604a3f16cf1d909bcf77a012802410fc1;
mem[513] = 144'h02f00f0208b4fbab00170ca4f9ea04ed0328;
mem[514] = 144'hfab5f8fef9e4080cf9d00208f852018d014a;
mem[515] = 144'h070bf06df904fbbdfbadf54a015505640a5d;
mem[516] = 144'h0ea007000e6d07a201b80bb400020f150fc6;
mem[517] = 144'h02ad002604370d4b0cd00c5c0aca0afdf706;
mem[518] = 144'h0a98f87d0d22f71109ed0d28f72f0ac4f382;
mem[519] = 144'h0d1cf21ff4b108050d42fda90b46028304e3;
mem[520] = 144'h0b3a0d2a0a94f5c60985f6c3f67b04d102d1;
mem[521] = 144'hfe670771fe840bbaf2cef7830f6ff561f2b2;
mem[522] = 144'h05d8f823078bf1b1f411fceb06f50dcaf328;
mem[523] = 144'h07be02aaf9c6077cfea1f050f9ee0ac6ff06;
mem[524] = 144'hf4e3fbe2feaafac60630078bf368f21df591;
mem[525] = 144'h0e6d01eafcc407cff7d10bba03f4026a03c1;
mem[526] = 144'hf8dc0a04064f05730afb0cf00dec0bb50a9c;
mem[527] = 144'hfdaafb0df9870f5e0409f3def0a1f575f70f;
mem[528] = 144'hf26af80f0c0c016af707fafc06d501d40c0d;
mem[529] = 144'hf1a409a6fe2000f802ec043709020357f14f;
mem[530] = 144'hf750034cf38009b80ee304450f05042e0b6f;
mem[531] = 144'h017e0957f252f57307030d9708cef7c0f409;
mem[532] = 144'h046b0b56ff1407cfff3d05d4f43a01100865;
mem[533] = 144'hf12ef6b9f0eafe040702f1e909ce02fcf331;
mem[534] = 144'h00d00f070b7f0328f3b5fffd0be1077e07ee;
mem[535] = 144'h0b120bbaf844f5f20350f41907de0b36fb4f;
mem[536] = 144'hff2d0f5d08f3fcfff2ee0f1cfcb10fa80a92;
mem[537] = 144'h0681f0b104f3fda0fa33fa510e8d0c5ef147;
mem[538] = 144'hf737f35d08b7f40afd85f5b6fe9af9eef673;
mem[539] = 144'hfad6fbc8ffb2f131fef50ed4fc19fb3bfed9;
mem[540] = 144'h0fcdfc22f16ef21a0747ff64f3a5f8b40b41;
mem[541] = 144'h00190bdc026d088f05d6041c08b302f20286;
mem[542] = 144'hf98e01d7fc19f22908f20bf0fe0f05db059d;
mem[543] = 144'h079af566ff4ff391f16d0844fc3d0f75fad9;
mem[544] = 144'hf0e80a370378020e048c00480a63f03ff50a;
mem[545] = 144'h071b0977fe9af2640a4af802007cf8920be6;
mem[546] = 144'h0a510883041ff0e20dc7fff0f5d0f306f63e;
mem[547] = 144'h091af612f61d0a39f3e8081a034af53e0040;
mem[548] = 144'hf6a9f9d80f99fce9f8870f460cb7f1ff0ee9;
mem[549] = 144'h0cb00ff30483fb25fe15f299f8d805a5f07f;
mem[550] = 144'hfb230888008af0affd19f15a07330c8f0ead;
mem[551] = 144'h0baa0beb03880a29f1460216f0d6027ff884;
mem[552] = 144'h0014feca0d720cbcfaedf96defee05d8f2ae;
mem[553] = 144'h06f0f010f3e3f94f033b0457023e0669f99f;
mem[554] = 144'hfa45f2de00befcb2fd0606a6ffbd0a680196;
mem[555] = 144'hf1f10fad01e9f73cf38103990c150e990e05;
mem[556] = 144'hf20700a6f8c00d82f09b033e03e803cb05ff;
mem[557] = 144'h0659f3c5fa0d07f604be08dd06aff2cc0813;
mem[558] = 144'hf6c205dffd9e0af1ff2e0ee8f59909200948;
mem[559] = 144'hf39b0a1bf1540d6cf4ba09fbf0ed08970ec5;
mem[560] = 144'hf8060093f20fff05f9cf08e7f83b0f8efd47;
mem[561] = 144'h0a0e0e0601bafb5bfc460797f770ff310328;
mem[562] = 144'hfb240b13f1f108f4fc18f1e8f999f7dcf4fa;
mem[563] = 144'hfe480e77fd5c02c9fdc10b69fa1d0b8e06e8;
mem[564] = 144'hfaa8f5040b4bf526f454f5eff79d02110dc1;
mem[565] = 144'hf59b0f09fa31006af58302bff9f50ee0008a;
mem[566] = 144'hf83a036300ed08fc096e0635fa3df7d00bbc;
mem[567] = 144'h08130c840e38f752f11cf4170b500e810c72;
mem[568] = 144'h05d10b40f6c7fc9a014b05f3049c030a02cb;
mem[569] = 144'hf603fd9e0165fde4fdb2fc7bfa57f2d00a93;
mem[570] = 144'hfb7d06eefb7500bff7800bb5f5b7f111018c;
mem[571] = 144'h046706cf0c95f591fc7a08e70ed3f585f514;
mem[572] = 144'h0fc3f6f5fee202ea02def079f3ebf88ff921;
mem[573] = 144'h0a2b0b6c075f076bfc5dff000d890f9ef443;
mem[574] = 144'hfda703c1f14dfa69fc7901470bbef599ff3c;
mem[575] = 144'hfff20ba9f39b0b1200edf678f833012dfccd;
mem[576] = 144'hfb73f08ff755f9d601d0f4caf5b1fb410501;
mem[577] = 144'hf39b0dd70bc404220835f3e8f455f790025c;
mem[578] = 144'hf54b0cdd059102270394007cfd100386f1ee;
mem[579] = 144'h0d2e0898f9520eb3f0670342fdd5fa4bf7bd;
mem[580] = 144'hfaf9f277f9e3f0b6f27cf6eaf225f74cf791;
mem[581] = 144'h0711058af33bf2dbfd19f107fc2d09bff834;
mem[582] = 144'hf54e0ace05a2f9630bdbf23909c40c0e0bf5;
mem[583] = 144'h035f042bfe4d0cc7f3d9f6c5fecdfaa8fbf3;
mem[584] = 144'hf8e3fab1fb5c02a4fe2cfbc6018e08150934;
mem[585] = 144'h0c49f372f40a02a80c89f1790d2004f5f026;
mem[586] = 144'h0a7ff71efac6f62ffa87fb130a140b4bfd08;
mem[587] = 144'h0dccf1b7f586ff76fd9cfe55f7fafc3f069a;
mem[588] = 144'hf6db0e98fc3106b7fdfbf6f306100b7106aa;
mem[589] = 144'hf9c60d4300d2fc650f470f0d042c047cfe79;
mem[590] = 144'hf30d0cc505cbf04efd08043b026301b70918;
mem[591] = 144'hfa160cf00d95f2ab05f00f38037afb2101af;
mem[592] = 144'h0c68f5b3049ef4be0c3301650a0808480036;
mem[593] = 144'hfb0a0aef025affe2070607d10c05f33af56a;
mem[594] = 144'hf0e6030fff40f26f01d8f1a7f75ef98a0512;
mem[595] = 144'hf2c409ff066effa8f22ff33d0ad2fa3200ce;
mem[596] = 144'h0ca207ec0e74f3620b17fa03fbaffe18f31e;
mem[597] = 144'hf3cbf271f26d0869f007f33ffd6107f9f0f8;
mem[598] = 144'h0311059405d7fb6bfb5400ddfe79f149f57c;
mem[599] = 144'hf669066af8f70e680b8dfef6ff8bfa220594;
mem[600] = 144'h0a40f2910623fa5bf326fc4d0d3b0231f1c3;
mem[601] = 144'hf79ef38afd3706bb00cb09390aa70d110b2c;
mem[602] = 144'hf998092e0cd4feed033bf940093d0cc7fc15;
mem[603] = 144'h08a9fe55fc07070af70dfdeb0cf109b20185;
mem[604] = 144'h0c3ff5dff9de07000279fbdcf30c0cc709a4;
mem[605] = 144'h0622f75e063e0feaf67607adfec1fb72f205;
mem[606] = 144'h0102f69709a8fc390ba90fb4f1a6f4d904df;
mem[607] = 144'hf2ab07180428f02c0f7307090f43013bf134;
mem[608] = 144'h053efad8fbc1fecffc39fc4f0c53f719f0f3;
mem[609] = 144'hf22df1a9fc6703110f37028df69e0e50f065;
mem[610] = 144'h0e90f1f8f98bf7df0a920afef63c0889f096;
mem[611] = 144'h0ff6fd7ef76ff7df067efe580409fccdfc39;
mem[612] = 144'h001e010df3a00dd2fac908100fa1f324fd1b;
mem[613] = 144'hff41f6c60cdafc550160fc95f209095307c9;
mem[614] = 144'h09dd0d54f5cbf48e09d503f8059cffa6f8f0;
mem[615] = 144'hf819fca5f05d000b00c4ff9c004f0767fa20;
mem[616] = 144'h0fcf0fac0d9ef8cb0390fc1e01060952f975;
mem[617] = 144'hf4f00317041af5980a690531f86c0743fab4;
mem[618] = 144'h0313f9f205550807ffc6f6d8fa5df607f9ab;
mem[619] = 144'h0c9b07d20955018cfbc10c79fbc4f9a3f7ae;
mem[620] = 144'hfaa7031c01adf1cbf93a065fffb4fefdf815;
mem[621] = 144'h00710e56fe61f0c40468049ff4f507dc07d3;
mem[622] = 144'h016ef210000306acfdd601200c3c0555013e;
mem[623] = 144'hfe6c017f01cdf8dbf1b1efd0f598f38e0744;
mem[624] = 144'h0642f3af01680af608d6f529f4dcfd780c5c;
mem[625] = 144'hf99cf2af054403f104e50d05fd0d0a640210;
mem[626] = 144'h05c3f6f70062f43d0e7a02dd0692f88bf919;
mem[627] = 144'h0748f9970e830583098304bef8b8086e09a6;
mem[628] = 144'h01fdfe83f3c003b20591fbc4f6c6f3dbf432;
mem[629] = 144'h07c4f175f816f4bb020e01120e4ef8c3013a;
mem[630] = 144'h0b240f15ff03fe44f3dc0ae8f935026e0b1d;
mem[631] = 144'hf04908eef330fa94f604f630fc66f4c309e5;
mem[632] = 144'h080ef8aefdd8fb7f049e01b7f4f60d5df1c7;
mem[633] = 144'hf132fbe000580c79008f03ab0d17f829fb7c;
mem[634] = 144'h008e0a74fa3afcf90a010d0cf98300770eff;
mem[635] = 144'h0699f30f0039f77efb44055cfcc7f28808b9;
mem[636] = 144'hfa1e0c26f24e082f09160172fd1802e8f73b;
mem[637] = 144'hff64f1f0fc3d08e8fef30ee6fdd2f054081d;
mem[638] = 144'h007f0d4cf5e8031b0ef2fea0f1e80fe0005c;
mem[639] = 144'hf7e6fc90f55bfbe00ed9f10e0ee90871f5ce;
mem[640] = 144'hfb08051407a505ca0d980d700beb00b4035f;
mem[641] = 144'hf37f0fadf57708d005e4023809fcfe2603a7;
mem[642] = 144'h0b870bb7066501d4f2520619f5c6f1410f25;
mem[643] = 144'h01dc05baf9ac0d280d12f1ce0076f53e0572;
mem[644] = 144'h09400949efd5043ef3560357f93009840805;
mem[645] = 144'h0112002dffc9fc17f1d8f6d7093afd270c2a;
mem[646] = 144'h0af7f1bf038e0ae8fae703d2075d0e4bfe96;
mem[647] = 144'hfaa2f8b30b9df627f284f39efc110fa4f2ab;
mem[648] = 144'h0dbd0387034a03fa025afa7cf5d70889f85d;
mem[649] = 144'h0357f61d0dd9fb1dfc71f26e0899f518fc95;
mem[650] = 144'h012f0bd10b630a90f78ffb600833f89d0a90;
mem[651] = 144'hf31bf90af67cf8cb0d54f1770c8e0aa8fe88;
mem[652] = 144'hf9d9fd43facd0f6af2a80e340cd00449f832;
mem[653] = 144'h063502230bfa0c8afdff01c009aef186f8b8;
mem[654] = 144'h00f5f3580b0ff4ae0660f0750cddf094f374;
mem[655] = 144'hf0e002ba0241ff3d08600c1f05e5fa7f0505;
mem[656] = 144'h0887f83401e20367fb36f522f8b9f6eefc6a;
mem[657] = 144'h0f2e0dc4f2210132075efc200705ff69ffa8;
mem[658] = 144'h0e0dfd3209e6013b0c3304b6009ff9490863;
mem[659] = 144'hf4920b56f4d303940cfbf0910c5c05e50f53;
mem[660] = 144'hfb3af6faf9b3f03002cbfc450019f826fb23;
mem[661] = 144'h04520e64fc48f8b8fc35fc1e04def89201c1;
mem[662] = 144'hf764f0ab0d780cadfe85f234074604020fbb;
mem[663] = 144'h07c9f3dcf480f262f8bb0585f662f893fabf;
mem[664] = 144'h06b70d6605d5fe08fde5f7f80fa7f872f98e;
mem[665] = 144'hfd770148036a0ccdf678f853fd3ff7e4053b;
mem[666] = 144'hfb9404950656fe6cfb5affa30445f4700875;
mem[667] = 144'hfa53fe69091ef2ab04bf059c0dda04b2f817;
mem[668] = 144'h06b0fa460fa4f98703010e71004ef7ca06b6;
mem[669] = 144'hffe5fdbb04c9f776fa2e05e10c18f8320257;
mem[670] = 144'h023e08970bb90b1d0be7f19f00c2fa17ffeb;
mem[671] = 144'hf5dafadbf275073c02f50f55fa21ff010108;
mem[672] = 144'hf61bff460d8206b20153fcac037dfb13fdc3;
mem[673] = 144'hfbe4061104aef2cff7c706c40391f7620441;
mem[674] = 144'h05c40528fa1bf23401ff03f3f97a01cdf7cc;
mem[675] = 144'h0acd0be501c6fa510425f946f59304960dfa;
mem[676] = 144'hf70bf9cefbd0f6e0f3ac019d042dfffffe64;
mem[677] = 144'h0ea3027bf86ff99300280d3d0f35f6e00eff;
mem[678] = 144'h004306b6f551fd8ffe92f99706a7ff1ef8fe;
mem[679] = 144'hf9020b84066ff53cf3380faff37af4d20006;
mem[680] = 144'h049af857096f053105b20bb109560e52ff50;
mem[681] = 144'h0c68fcfa0fd902580716033f0a530547f46f;
mem[682] = 144'h00450c910d6c0d34fec1f736fcbdf990f58c;
mem[683] = 144'h02140c090b9f0d18f1f20ff80d430e5a0f8d;
mem[684] = 144'h053cf911fb4ff253feca05980581ffdb0af3;
mem[685] = 144'h04a604abffd7f0e505f60ead0d170fbd0524;
mem[686] = 144'h01bffef6056008b9f4eb070bfd62fe49f9ad;
mem[687] = 144'h05bcfe43f8c402370395f907f416045108f4;
mem[688] = 144'hf29c0f69fcc402cc0210f4c4005701b00516;
mem[689] = 144'hfbd9089efd65f7fd0fb0fe140b93003c0e42;
mem[690] = 144'h0d5a08def9bb0f65f5fc0e78fece0f0005c9;
mem[691] = 144'h07340cae0940ff94f4130db10a3d0a44026a;
mem[692] = 144'h0a51075cf3b2f273f7f7fc54fc8f00a1f629;
mem[693] = 144'hf7c6fe0cf82ff0220b8ffb5bf42ef90d07dc;
mem[694] = 144'h0564046c0b6ff86bfc160c07f6aff3d7fb4f;
mem[695] = 144'hefe50f6e0478040b0c6304cc06a607abf3fb;
mem[696] = 144'h0d85fb030b7eff26f5e5f251fd0a0b920723;
mem[697] = 144'h019f0c220e7ffe39fb740e4afc1aff19fc59;
mem[698] = 144'h008403880364f2f307a706320d970b6ef085;
mem[699] = 144'hf6fa0ab1f134fc53efc9f4b7f5abf6dc06ed;
mem[700] = 144'h06edfb9eff1c025cfee40090f6a604b0f3b0;
mem[701] = 144'h0adb09500a760e19f7eafa290c4e071df3da;
mem[702] = 144'h0e99f829f2b001daf9aa002ffc7104fbfe0b;
mem[703] = 144'h00e0fa43f8e00455f60305d50727fc4afdc0;
mem[704] = 144'hf1690b1ff416fdeaf7d0074b02aa0459fa96;
mem[705] = 144'h075600f6fd0706a00e0909a30ac60a7af042;
mem[706] = 144'hf836f7d3fae1f7e7f712f5a80d9b060cf467;
mem[707] = 144'hfd5b0ae9fe0efce2f1df006ef5ccfc1cf27f;
mem[708] = 144'hf26bfea406b2f52afd40054b05bff08a078d;
mem[709] = 144'h041f03430646f76e07c00148007e05c20e2a;
mem[710] = 144'hf2d8fec7f888064cf1c7076af570f8c00764;
mem[711] = 144'hf0c504bcf68608320b7ff707f081f51f0ead;
mem[712] = 144'h083e086bfe0dfc2f0cd80b97f71702a4fc89;
mem[713] = 144'hfb6dfa3703e8ff1a0186f74e00cbff65f9f5;
mem[714] = 144'h0618f1ddf9f40d3e053809e50f710b65f561;
mem[715] = 144'h01620241fcb50c8c0ddf049ef47f02ddf99d;
mem[716] = 144'hf33f08cc00b80e690c26f56e00eaf0160666;
mem[717] = 144'h04d00a660827fe36f408088b055cefdb0889;
mem[718] = 144'h082e04abfa0c0af40a89015d0d390acf0d2d;
mem[719] = 144'h0a6e0e4ff34afb34fc98faf00ee5f30907be;
mem[720] = 144'hf08103c3f3e600dbffbb0fa10bebfdfcf9fa;
mem[721] = 144'hffab087c072c060d01930ce8ff49f1def3eb;
mem[722] = 144'h0c5601bd0545fa180676ff21f6d006c80427;
mem[723] = 144'hf8bdff6b0fc6f2a508b90bccf315f380fd22;
mem[724] = 144'hf2a1fcf60ea3f2f006e5f078f4290c10f681;
mem[725] = 144'h07e0f6ddf1d0fec707def5c20104fde90799;
mem[726] = 144'h015501bb026805ccfd7c02b300f008890179;
mem[727] = 144'h0620f19afc44ff87f9360a7e0fec098dfd13;
mem[728] = 144'hf50e00ad0705fbfd0f930ac0fc54f4c500ad;
mem[729] = 144'hfbf1fbd8f7d607920478f5aff16cf9300a64;
mem[730] = 144'h0f9a071a003003d7f32c0194057ff463fdf9;
mem[731] = 144'hf58e08fcf36607be0d82fd910b7ef27506dc;
mem[732] = 144'h0666f96d0ba00f760805f0f4006800c5f4f8;
mem[733] = 144'hfef5099e0fa1f365f54d045d06acfe56f065;
mem[734] = 144'h04e2fd8807240a46f951f0260974f8f30e59;
mem[735] = 144'hf8ce0f35f59907b0f40e004e088406b2f3e5;
mem[736] = 144'hf06cfab703a706170000f08afe1cf5eaf171;
mem[737] = 144'hf6990bacfc51f7270d9c07ddff060d760f1a;
mem[738] = 144'h0d6ff73b0b75f99d03170af4f00801cc0b64;
mem[739] = 144'hfa11ff85fdc702c807b0fc19f1000b78f5c4;
mem[740] = 144'hf9e9f80dfa50f44a0bd40a05f23cfeb90894;
mem[741] = 144'h0b4705840936f4600af1fae9f43801b0f835;
mem[742] = 144'hf972f2cbf3c208a70f820412069c07da020f;
mem[743] = 144'hf8890a610959f889f3d5fbbdf24108390ed9;
mem[744] = 144'h0b08fb3608c50e8f0e17feedfda107a5f3c1;
mem[745] = 144'h010dfe0afdb5029a07e7fc920f800512f338;
mem[746] = 144'h077f093c0b60fa45f31ff844ff27f95ff43c;
mem[747] = 144'h064e03d80f0e0e8ff1e1fae6fdbf0a5f044d;
mem[748] = 144'hf2730cf90021f2d1f1a5f123019309b606a6;
mem[749] = 144'hf84ef1730375faa7f095f0b207d0fb7509dd;
mem[750] = 144'hfb65f9e2045008a90a510347094c032202c1;
mem[751] = 144'h0f18fb71fc80f518f8020628fca1f74903ef;
mem[752] = 144'hfbebfe97feebf62003690ceafb56fbfafa47;
mem[753] = 144'hf1ed07a6fa75f4ec0b0803d5060e0845f692;
mem[754] = 144'hf99af0380860f15802c2ffe70d0201110ccb;
mem[755] = 144'h029df217f9bd0c2004070c4df05306d20fdc;
mem[756] = 144'h0b600298093ff24c0a17fb32f1730f5bf7b8;
mem[757] = 144'h0577fa5df95afc06f7960b3d049cf66cf2cc;
mem[758] = 144'hfc380a3c008efca709df0850f008f094f259;
mem[759] = 144'hf3280d6d08bb03e3076f0651fc8df2c70463;
mem[760] = 144'h0f67fb69fefef533fa4008b0f25702c1051f;
mem[761] = 144'hf1fcf38cfd620741fe6ffd9cff3700630e09;
mem[762] = 144'h06a7f852f040f7530525f75bf38b0bd40973;
mem[763] = 144'h09cffaf7fa380a43fe620fea0f2c079e0a95;
mem[764] = 144'h0c84f82a0e49fb1004700c52f476f97bf136;
mem[765] = 144'h0949f6eff474085cf413f2edf825015a030e;
mem[766] = 144'hf857f384fb47f7340c740da9f823fa25fad8;
mem[767] = 144'h0129f6d1fb3e0cc9f712fac20c530e20f995;
mem[768] = 144'h08ccfa6f01f105fafa3ffaf8f8cdfcdef89c;
mem[769] = 144'h008d0d5e025d04e2f1def4d50840f6c508f3;
mem[770] = 144'hf25908880c0600e40efd086505c20c05fb25;
mem[771] = 144'h060ffe9ff7e301b40754011c0ef5026600a7;
mem[772] = 144'hff2d09dd057cf89af77006e501b9023903a3;
mem[773] = 144'h0f00044a0adcfe7bfacd0edbfd08038405f2;
mem[774] = 144'h0115fbfdf296f0c90196f7eaf61c0b26f2a9;
mem[775] = 144'hfc34f2be09030ae1f7ba04a3faa00f72febd;
mem[776] = 144'hff9408aa03e0ff4bf280085409d80832fd97;
mem[777] = 144'h035100fa0d0bfc8df0aa033f0db60403fd32;
mem[778] = 144'h0407fd3802cbff7405cbf8610f1501340732;
mem[779] = 144'hf4d0f1ca056ffa35fe73fff60ae8fb8c0b4e;
mem[780] = 144'h0634026a0e3bffa40945f76f0c3ff2a20cc0;
mem[781] = 144'hf476f55904eafc35f6eb08edffbbf16b0f70;
mem[782] = 144'h0eb7f462fffa04a5f46d04e006d8f4f40994;
mem[783] = 144'hf1550342f9c1f730fce7fd9b078ff88c0dd7;
mem[784] = 144'hfad8f8c8026c0975fe4e0b8cf5faf8830291;
mem[785] = 144'h05a3f1b9ffe607a1015cf603f10008350b6d;
mem[786] = 144'h088ef0b20be1f831029df5c1007afc94ff8f;
mem[787] = 144'h0ba4030e0ebff995f67f0c900c6a07b70c54;
mem[788] = 144'hfa60f19df381f148fb150eaf0c810bfafb10;
mem[789] = 144'hf017fb60ff8200db0eda012c0622093c09ed;
mem[790] = 144'hfda60d30fbd60eb209ccf6ff078d0cdff64e;
mem[791] = 144'h04440da30050f657f237f0cf04ea058af80c;
mem[792] = 144'h0dd8f36005fe0eebf06af586f2bbf2030b71;
mem[793] = 144'hf38bf474f40f0c5bf64af2ec05ceff4808e7;
mem[794] = 144'hfe3b0e130b29f304055503d0fedff649f2d6;
mem[795] = 144'h0613089c0087f42803ba093dfc9df5350746;
mem[796] = 144'hfdf7f2d606760ca9f2b1f18cf3f2064ff797;
mem[797] = 144'h086bfaa5075102ed0477f0eb0e870e78f6d8;
mem[798] = 144'h07b1f49d0785f1f0067205d3fc1609eb0038;
mem[799] = 144'hf60e0cf2f04a0a180094056dfc6d0dea0659;
mem[800] = 144'h0722ffd1f3c1f077018f0eb60ccb0773f7ae;
mem[801] = 144'h01c90db4f4d9001dfc8afe8af5320fb4f60a;
mem[802] = 144'hf2b7fc90f54ffce7f331062100b4fea505be;
mem[803] = 144'hf6bff37ef7020c8d095bf346f197081b0492;
mem[804] = 144'hfeb8f4b5072207cf0ebd003c02baf7b1071a;
mem[805] = 144'hf28ff4e1f748016af4650c64063ff1f5f49a;
mem[806] = 144'hf76b0aad0557fee6fe5df8f50fbc056b0c77;
mem[807] = 144'hfab00c31f80008fffb1ff94eff8ff8eef576;
mem[808] = 144'h00f7f257f5160d7806bf0ec20c8afd010e75;
mem[809] = 144'hf5a704890f470e7ff8130e3efe54fa76fdab;
mem[810] = 144'hfdb0fb67f4a70d52feb7f2da055c0af0f23d;
mem[811] = 144'h05fefbe20f6608a3f60afb92f7f20b42fc70;
mem[812] = 144'h04fd0053f61dfeca0e46f4e0f522083e0154;
mem[813] = 144'h08820621fe700005fe05f3b3fc760475fdd4;
mem[814] = 144'hf4d705f4006b0c95f4c1ff8303c2f6f5f761;
mem[815] = 144'h06950b30092703610ca7021c0a5f023afd2b;
mem[816] = 144'hf804f8b0fcfaff17015701eb0512f9bff017;
mem[817] = 144'hfc680c46f879f2cb054b072e056504b1fda8;
mem[818] = 144'h0752f8140b350e52f5540d42f34bf6a90688;
mem[819] = 144'h0037fb00fca8096a0f2ff6c9057201c3feeb;
mem[820] = 144'h0592ffb90c3e0e3cf9a405510102f3c3f3c0;
mem[821] = 144'h022af2b4f70efaa2f35007fdf9a80fa5fa0a;
mem[822] = 144'hf0e802f9f0d70c5002ca08e1f64ef14c058d;
mem[823] = 144'h0430f7c30331013afd890cfaf0bff89f02d9;
mem[824] = 144'h06650eaaf8a4f06d0ccd0c2d0c240c7af7d2;
mem[825] = 144'h003f0ea4f72c027f0085f600f2f50c97f60c;
mem[826] = 144'hff9df20afabbfcd20e45fa0af14bfa4af0a4;
mem[827] = 144'hfd81f340f7c80e050a5808f3fe54f100f229;
mem[828] = 144'h0e560eb2f05d0db80918fb79fd54f2200999;
mem[829] = 144'hf2b4fda5f82e0955f85af232f998fccafecf;
mem[830] = 144'hf791042609e3f951f34ef0d0fab8f32c0829;
mem[831] = 144'h05c7f29d02f9fc60fa67f37307930a40fa3f;
mem[832] = 144'h029e0b49fdac0fa7f806f443fdf6ff5cf400;
mem[833] = 144'h00a4fd0ef773fc530f3009a5fa9cfc65f818;
mem[834] = 144'hfe55f6880eb40d6af344f5340fe6083bfebf;
mem[835] = 144'hfd9af873f72f08cffd6d06720f4009a1f30c;
mem[836] = 144'h025e0c88f004f715f4effdbe049bf4d8f5c9;
mem[837] = 144'hfacc07a4fa0ef6e00d12f4760aa003e3ff90;
mem[838] = 144'hf0d5f30e04cb0ba80fdcfd53f773ffd50360;
mem[839] = 144'h04e6fccb0210004affe20510f14d0032f511;
mem[840] = 144'h05e60d11001ef0a1042e033ef3800c04082d;
mem[841] = 144'h001f05410725fa62f7f10f1f0f5afb8df285;
mem[842] = 144'hfe5008baf6a4fe2d0416f8cd044a0c52fec5;
mem[843] = 144'hf99203bb085cf02a025ff60cfd00ffacf542;
mem[844] = 144'h08acf64b0d67f0d1f7420792fff30e930cda;
mem[845] = 144'hf66603400c0206220b83fbec095cffc0fc32;
mem[846] = 144'h00b30ec4033200a40e9cf224008809dd0e37;
mem[847] = 144'h0918f6e6fda9fd14fd5208ef04d304a6f7d6;
mem[848] = 144'h0da7f927f445fe6d0b0e0264f157f365ffea;
mem[849] = 144'hf0870c24ff8f0539f6e4f0e0fdd8fca4fd2a;
mem[850] = 144'h04d7052a089ef3def4a6fdb2fb7c017afba7;
mem[851] = 144'hf7ab0286f897031df7cafb8af70c056a0eeb;
mem[852] = 144'h0af8fa04f343033707d20b2ffd0af1e7f634;
mem[853] = 144'h036c0acb0fc8f4c5f39bf00e08a70f1c0657;
mem[854] = 144'hf8baf7810c6e0b630746f35afaa205c5f174;
mem[855] = 144'h0d3ef33efb4f01ca0727f99ffcdb0230fcb7;
mem[856] = 144'h0ebdfbc9f67cfde2f8a1f0a4f2350df80eed;
mem[857] = 144'hfd04095f0b3ef1420445fb5df93701430ced;
mem[858] = 144'h03d1f5df0025f213f0acff2306bb015cf405;
mem[859] = 144'hf4a5f7d905130d68034df9850c87f6d50f7e;
mem[860] = 144'h0c300b4cffdef1ebfc020a6f0ad803990bd3;
mem[861] = 144'hf9ca0e9d0604079bf224f3e7f5fb028cfc64;
mem[862] = 144'hf4ee0318f06902e4f027081b0b1ff0780932;
mem[863] = 144'hf08ff2d0049a0f180692fe0cf80bf60ff6b8;
mem[864] = 144'h0193f66bf1e50499ff8dff88f551f58a06b8;
mem[865] = 144'hffd208e903bb02a4f8d5f89b043e0cf60771;
mem[866] = 144'hf56c0d450c0002f1057df1560401fb6ef8f7;
mem[867] = 144'h083dfdeefd6301d4ff5df00bf2b0011f03d7;
mem[868] = 144'hf26df90cfbdafdf4f90d04eff85df668fb89;
mem[869] = 144'hf3fbfbc2f60d01ef07d109510f940b590313;
mem[870] = 144'h0639f0befe68fc21feeffd41f472f12e0044;
mem[871] = 144'h06fb0e9af527fa350d800296ff03f623046b;
mem[872] = 144'h06ddf31ffe7af1aef619f5d1fe01fabc05ff;
mem[873] = 144'h043efd90f94efcb0062f0f45fa2ef5e7fb97;
mem[874] = 144'h0ba30d2b09da0124f08ef219ffd7ff200801;
mem[875] = 144'hff190f6ef1460d07f4eb03b2f821f86bf7b3;
mem[876] = 144'hfaf901e2f785f60b0b8305330e49ff600322;
mem[877] = 144'h0149fe39f9340ebd010ef157f5b90703f86a;
mem[878] = 144'h0b5d089af7faf566f688f156013b079e07ae;
mem[879] = 144'hfe00ffbc0c9ff98c0b2df594faa3f7be0075;
mem[880] = 144'h0b090159044c097e09c5f0b303f2061c0754;
mem[881] = 144'h0e080ee7fde0073a0f42ff05f02602db054c;
mem[882] = 144'h0101f016f202fb800479f739fc950664f26c;
mem[883] = 144'h0957fd1a0fb9f9650546fc4cfb7b05edf4f8;
mem[884] = 144'hf850f2120d45f58dfa850022037d0bc8fcf0;
mem[885] = 144'h029cf40f0b2afa6f06f8005f0381f108f183;
mem[886] = 144'hfa5bf4b50b84fbcd03850d29faa0f7ccf968;
mem[887] = 144'hf378f57b00b5fd220617fbb10e5a02be0632;
mem[888] = 144'h07a9fba309a50b660f61f97d0c3bf2c502ea;
mem[889] = 144'h082af4a30e8f074c0828f45402d90ea30be3;
mem[890] = 144'h052e0070f0810183f19308ff080df2ad0495;
mem[891] = 144'hf99a0d12eff4f9cffdc8f74df7caf1810da2;
mem[892] = 144'hf9cdfecef705f41c081506bb082bf0cffa05;
mem[893] = 144'h0d15f816061502630ca702e5f63605c0fe23;
mem[894] = 144'h06d7fc5df2980a27f527041a0d1afe210bde;
mem[895] = 144'h0a12f0f1f7f8f015f64001ef00a8f53904b1;
mem[896] = 144'h0c6ef660093f0576fc24fed706f1f0bf08e2;
mem[897] = 144'hf90a00230b4bf98bf8bafa5fffb60d88f02a;
mem[898] = 144'h044707c7049206fafbe80551f03ef37cfe39;
mem[899] = 144'hfc58f1a30d01015b0b25fa3107760e8ffcbc;
mem[900] = 144'h05fcf1e90ff6f63bf00afbca043e08aaf738;
mem[901] = 144'h0bc6f2580aec04cff3baf734fbadfe070ed9;
mem[902] = 144'h07ef0bf407c80375f3e601e10211f9f2f77a;
mem[903] = 144'h05c00038f4f30cf1097bf54cf90dfda0fe1b;
mem[904] = 144'hf8f405f005620a30fd0d014b0261ffa9fee9;
mem[905] = 144'h0474ff5bfc41033ef82bf7e00ce00b380090;
mem[906] = 144'h053f06e10eaaf8250875f904fb5ff35309de;
mem[907] = 144'h041bfea9f3feff3bfa55ffe50631f046f320;
mem[908] = 144'h001fffd7088df58dfaf9f90f01f80863f177;
mem[909] = 144'hfbaefcf5020c0ea401a10f6203390957fd08;
mem[910] = 144'h02fa0788f7e4fbd10c380cf00bbe084902bb;
mem[911] = 144'hfd19fdd0fc65fb610afe0d91f87e09f5f1f0;
mem[912] = 144'h0cb9f03af2e0fc68f5d400e5f06bf2670bbc;
mem[913] = 144'h065bfd76f4be0f3dff6c0f03fc39f7460673;
mem[914] = 144'hf0720992fa250083f4ff0bcd0170f033f54a;
mem[915] = 144'hfa2cf84a016d0f7d0dfffc5d034204130c3a;
mem[916] = 144'hfdd6026af543f5ef020905ec08450db70530;
mem[917] = 144'hf42e0c8c00e409320f460647f4d1fa550239;
mem[918] = 144'h0973f3aefe1404d10c4d092cfebdf542087f;
mem[919] = 144'hf762fd4c0cc00b9c0ac4f12104d6f3d5f89c;
mem[920] = 144'h0bc20d33f83dff2203b006610f10f2cdf3bc;
mem[921] = 144'h07850a53037f06d3f601f5a1fb60f698fd40;
mem[922] = 144'h041e0d30fade0cd8029c0db402230af4ffd4;
mem[923] = 144'hf184f2defd5a027406510316ff3007e90e33;
mem[924] = 144'h00620b11fd2bfbf6097a015702130d9cfce2;
mem[925] = 144'h0a7f0a850cb60fa20ba50d9bf4e8f95702e4;
mem[926] = 144'hfbd50ea10816fb4ff97406b7fe620ab400ab;
mem[927] = 144'h00bffebb010a0888fe830e2bfb200a31f7b5;
mem[928] = 144'h011bfc06fd3c023e008100720636028d09e7;
mem[929] = 144'hfd79044a0dc9f00908a0f1a500e2fdaff764;
mem[930] = 144'hff070cd0044cf855fc74fb0600480316fcbc;
mem[931] = 144'hff5ff79f02dbff40f414f5c8fe700a34013c;
mem[932] = 144'hfa510ac1f5840dc0fe36f32cf778f2930ea1;
mem[933] = 144'hfba3f77d053a09dff69304c90f06f4b90239;
mem[934] = 144'hf18c0b4c032af92df542f9d70c83fea50c5d;
mem[935] = 144'h0c11044906680d84f17f0f5e0541f4e2f1e9;
mem[936] = 144'hf3bb01c0f08404da0d95f117022e0ba6fee3;
mem[937] = 144'hfbaaf9c408e0f8030ad5fd21f8a900520c54;
mem[938] = 144'hf2b10d6f028cf028fd430d4900070c5b0f64;
mem[939] = 144'hf06d09bb0f3df7d80e43f0a0f33103c1f0ad;
mem[940] = 144'h026cf2f10899fe9b031406dfff91f51ef3fd;
mem[941] = 144'hf874002ef267f88fff2bf84f0af108f2febb;
mem[942] = 144'h00d6fbc0fdeeff340d2709e0fd84050df59b;
mem[943] = 144'h06080f600c54fe3cf2b8f913064a02220a06;
mem[944] = 144'h0a010aa9f5bef04df59a0cbf0cb8fca9f6f3;
mem[945] = 144'h00830d15fac10ee1f922f032061bff9c0460;
mem[946] = 144'h0c5c0f240bf5ffc1095ef0d2f7de04e20d39;
mem[947] = 144'hf8e60693f24f05af0611f68b0d2ef5d70133;
mem[948] = 144'hf178fb13f34affabf526f186f924f205fdd0;
mem[949] = 144'hf2d9088cfbc805c4f7e00b8b06990bda023d;
mem[950] = 144'hf02c0b7c062df30ff6e1f2d4f3890d1df164;
mem[951] = 144'h03eb01430da601ce0b2c0283f016f6be0084;
mem[952] = 144'hfc6c02cf03e9f80b0417fb84f9ecf33005b5;
mem[953] = 144'hfc7f0c95f9bff192f6acff65ffc4f17efbf7;
mem[954] = 144'hffccfbd5f92b06fa09ea023508c4ff53fc55;
mem[955] = 144'h0cf2004e0bbafdc8ff20f86bff3200e205eb;
mem[956] = 144'hf98d076cf7c0071ff30b0d79fbdb0da9f5a7;
mem[957] = 144'h0eba0d9bf4cb026706cef75a0226f945f0f3;
mem[958] = 144'hf8f9efe1014bf1220f8b0ec0fdcd0261ff55;
mem[959] = 144'h03a10f0df7e802f70e9df6fc0e97fcb30f50;
mem[960] = 144'h0b6606110f93fc07f226f4d306c3fce0f7d1;
mem[961] = 144'h0648fa3b005af4b10b10f29f08e3fb90fb5a;
mem[962] = 144'hf3a5f3cefbe80b5cfcca0cf8f171028e005b;
mem[963] = 144'hf50c050c0265ff51f28802fcf01a0809fe1b;
mem[964] = 144'hf9ecfb230364097b06820bd1f0b60f4409b8;
mem[965] = 144'hf5d8ff96fa15f8faff83fb1c0884fb3c0321;
mem[966] = 144'h07420c91f756f0860401f283f35af17501a5;
mem[967] = 144'hf1c9f42000d6f5f5fce103c006dff95401be;
mem[968] = 144'h08acfb1a05710590f4df024909bf0460fd4a;
mem[969] = 144'h024b01200f00083206f80959015ffd31fba3;
mem[970] = 144'hfcca034cf40a0b5d0a350f6004fbff79ffed;
mem[971] = 144'hf9d509bf01db036400ee065d0b450a47f858;
mem[972] = 144'hf7a8f556097d0ae60799034ef28df9110a3b;
mem[973] = 144'h0c9804e30808f2e6016d0de407cf0decf4c8;
mem[974] = 144'h0bc2f2c2099dfe30f123fd99f83002e0faf2;
mem[975] = 144'hff50f7dc092bf06ef65d01530769f250f45f;
mem[976] = 144'h0092f00cf84d09760f400b3ffb4c06bfffc0;
mem[977] = 144'h00a9fae40f0103070e3d091ef1ef04cdfdc9;
mem[978] = 144'hfe29009b0889072e0817ff120aef0d1e0d40;
mem[979] = 144'hfca7f3d00cbd07e3f34f03030052f717f5e1;
mem[980] = 144'hfda6f154fd2ef5e9016804dcf95300b1098a;
mem[981] = 144'h039b097c09ee00a9f95efa8ef5acfccbf45a;
mem[982] = 144'h0542f05ffe87f4c1ffcd01cefc8af905f4d7;
mem[983] = 144'h0660ffd4f8c205a00200f8f4ff1108ea09d3;
mem[984] = 144'h0ab1fa35fcd4f881f767fac0ff49fac5fb39;
mem[985] = 144'hf2d8f21b09fc09250320025f0fd4faabf6fd;
mem[986] = 144'hf87d0347f00e00bcfe34f8500844f1d5fbd6;
mem[987] = 144'hfe47f0d404d4ff3af5e3ff67feb1f83af691;
mem[988] = 144'h06edf5aefee7f461f04efd62030ef80df00c;
mem[989] = 144'h0d58f5720480f345f7d30d3a03dff3dcff3e;
mem[990] = 144'h0064f39a0137f808f89f0956f064fa5d0574;
mem[991] = 144'h0212035b0d9e072ffa34f94cf7130ab40593;
mem[992] = 144'h0641f8b8fde4f842f7b5f662f54ef114f73e;
mem[993] = 144'h02470f66fa91f3e6030ff4b30ce9f6e90a71;
mem[994] = 144'h051a0a3bf537f624f9640d21f17d0448f2e5;
mem[995] = 144'hf91df40efeb3f699f418f57af48ffd44f7e6;
mem[996] = 144'h03aefc7bf814f747f8250387fb5009320fb7;
mem[997] = 144'h0da6f9def331016f06b1f944f7aa0cfcf10b;
mem[998] = 144'h02aa095cf151fa5ffe8afb6206380a010f6c;
mem[999] = 144'hfd8bffc6f726fb33f02f0ca5f295fa20033b;
mem[1000] = 144'h002af05b0c1e0b4b0dd7f7f703f0f9f8f643;
mem[1001] = 144'h0a5cf5530e33f27af492fefd067cfae10c30;
mem[1002] = 144'h0ceff975f5ac02c40f51fc0c0946f1e2f80a;
mem[1003] = 144'hfc4f04bdfd3eff020ec800a20eaf094b0cf8;
mem[1004] = 144'h0885fa70f33d0e510dcdf1b70249f7eaf159;
mem[1005] = 144'h07c5fd570ee807f208f90fed0a350b5d07fe;
mem[1006] = 144'hf3a8f00a0f14f84cf06b09870d79f70f0235;
mem[1007] = 144'hfd0c0963fabcf830076909e70c07f575fbfa;
mem[1008] = 144'hfe30fb8209d70c2ef7e9fb4e0bc7f5adf825;
mem[1009] = 144'hff7a03480fbdf010050afb3803080a79f4ff;
mem[1010] = 144'hf96e0462008df4ec047afa7efa1f00d00fc2;
mem[1011] = 144'hf7c7f27efc99f7c7004f0dc400260948f91d;
mem[1012] = 144'hf7c60bb8f6740b31fc94fd8004c9f9e7f6c7;
mem[1013] = 144'h079f0046f6ceff68023cf03c0cf1fcbdfd05;
mem[1014] = 144'h0d68f5ac0357f0dbf31809930c580c5c009b;
mem[1015] = 144'hf753fd85f9e3f5c40921fe0dfe640234002c;
mem[1016] = 144'h0febfd39ff54fde3ffb901f2f6b20b20f60a;
mem[1017] = 144'hf1e5f219fd830866022800ff0880f18cfc80;
mem[1018] = 144'h09a3fc24f874ffa501de08f9f085f609f9d9;
mem[1019] = 144'hf793fb2ff4bb0a5f01a90e46f8030631f912;
mem[1020] = 144'h0951f6b20b060595f7530e8df647f5bb0893;
mem[1021] = 144'h0a67f3890767f551ff63054b035b06a6f06e;
mem[1022] = 144'hf42bf63cf65efdd5f6fcf008078bfafb0365;
mem[1023] = 144'hf6aaf7c8f695f87cf0c8079bf5ebff24f6ae;
mem[1024] = 144'h0e69fd8cfd27f8ab0a93f15df4ec0cf1f797;
mem[1025] = 144'hfb950c67f0c3f6abf897fa9106bbf463fac5;
mem[1026] = 144'h0e690e6e03f2fbda0c51061d0910f817f2e5;
mem[1027] = 144'h048f0753f321f2f2ff42f19b022efca800c0;
mem[1028] = 144'h0b07f0cef601ffd1f7d3001e036ef3cafa87;
mem[1029] = 144'hf02a09d3fe48f48e06c1f8e00778fefef88c;
mem[1030] = 144'hf52af0d1f05f076ff2d3f158f14309150100;
mem[1031] = 144'h053d0351fbb3fd3bff85f7c4fbd303fa0158;
mem[1032] = 144'h053f0dafff600cc5ff8809c9f1240200f69e;
mem[1033] = 144'h02e10a4cfbd708f4fcdbf14806a3f75df45d;
mem[1034] = 144'hf433f8d6f3c0f1c90dd40eed0742fb3209a9;
mem[1035] = 144'h0d2d0cb108c2fbd10fc103fe0ed7f026f877;
mem[1036] = 144'h0735f05501da013c04a2fbc103b50a06f9a4;
mem[1037] = 144'hfea1f24bf1c8f5f6005d01cb06ad089b095e;
mem[1038] = 144'h08c00d910d6f07450b1eff5a0014fb3df7e5;
mem[1039] = 144'hf35afe69fc20040b05bb0f430bea04ff040c;
mem[1040] = 144'hfb33067ffe73f06c0b41f4ce0a2b02adf29c;
mem[1041] = 144'h0f03fb4a0acf00e8f1780957f449f2500840;
mem[1042] = 144'h06360e4206d30b5df699f08d0f1cf1a2fa03;
mem[1043] = 144'h0e9e01c804dc06a7fe39f671048bf16f01e8;
mem[1044] = 144'h0c3df5780c240f7a02a4f53f0830ff850832;
mem[1045] = 144'hfe820801fc41fac9f2fc0b520bfc0c6f0608;
mem[1046] = 144'h0f18f53503f1fe030cc70403f957f0b606c5;
mem[1047] = 144'h02d7f2b50fcf099cfa9cf14a0e20fa92fe48;
mem[1048] = 144'hf303fa7c0cda0d1700e20dc1f2eaff5df3a2;
mem[1049] = 144'h018bf8ca04ad0933faa2fea606e3f68b0a16;
mem[1050] = 144'hf5bffee0079b0470f9b4052104140ddffa68;
mem[1051] = 144'h069b0b0606d0087afc270c71005c0e630028;
mem[1052] = 144'hf18905640c220dd30450f3c5faa8010703a1;
mem[1053] = 144'h04b5fe8e02baf57f0dbf0b330eb7f2bdf875;
mem[1054] = 144'h0eb1f677f34dfce5021df07ef0c0f33403f7;
mem[1055] = 144'hfe02fb50f8e302000b3401d5f697f269fa87;
mem[1056] = 144'h0f74fc29fc31fc5cf109f75e04c0fdd7f3a0;
mem[1057] = 144'h0986fbd80c2efdb30bcb0abf0394f37706d7;
mem[1058] = 144'hf69e0eb3f99405e9ff5f006502c30756091c;
mem[1059] = 144'hf5f30a780f810b3809870043f69ff66efd43;
mem[1060] = 144'h0dac0a8e0434f582f1b0f2fb0c4cfd490837;
mem[1061] = 144'h01b10b8a088d0b76f9fef4cff85705c40f4d;
mem[1062] = 144'hf6cc014ef5fdfcbafcb9fad70e5cf25309fb;
mem[1063] = 144'h082af6e4f4e5f80a00c4f3d7f7d50fb6f873;
mem[1064] = 144'h0607f972f9d70c970ca90ab30315042103e5;
mem[1065] = 144'h0d1409a60c0509d7018506f0069af651fe7d;
mem[1066] = 144'hf002f90c09a9fa270b10f2ef0a9f027fff90;
mem[1067] = 144'hf429f48df6c7f7a2f0600c730c85fc8e0278;
mem[1068] = 144'hf8eeff7bf52afd7303f9055ffab80565f3d5;
mem[1069] = 144'hfb26f1db0b8f0227fc0c074c076dfc0efe12;
mem[1070] = 144'h0518ffcff406f6e4f4fd07960827fc57fff7;
mem[1071] = 144'h04ad0b16058bf449f6260fa7004ff9790587;
mem[1072] = 144'h02330c8008720115fe5609d604ebf3c30d31;
mem[1073] = 144'hf514fe4bff500ad3f7ae0575096d01a2f12e;
mem[1074] = 144'h01c0f227f870044bf39cfa9e08e5f5410346;
mem[1075] = 144'h0d1af36505b2093f00ed084bfae2f15f0cfb;
mem[1076] = 144'h0201f06903ea0e67034505ee0ca70d4e0ec2;
mem[1077] = 144'hfb8a01b4ff2cf7e50db201ad0b42051ef7e6;
mem[1078] = 144'hf1390896002ff2f2f0c1f03108590d6e0beb;
mem[1079] = 144'hfa6efb910a9b05400977ffe2095b06d50a83;
mem[1080] = 144'h0370f462f8e80095ff750cfe0455f8290ed1;
mem[1081] = 144'hf6def3fd0a1102f00b5c03160b520671f847;
mem[1082] = 144'h0e4e0a8701150fc7004308faf53ef1c80ee8;
mem[1083] = 144'h07adf80dfe510994fdf6009908d1f146f0ef;
mem[1084] = 144'h04c0fd520d5b0446f574f657fc97f4a50bc9;
mem[1085] = 144'hf13403e5fd120188f4faf7bffc68ff6bf609;
mem[1086] = 144'hfd52ff4203e4fbbcf659f94ef9cff3ed02a4;
mem[1087] = 144'h03750ca6f43b0c7ff13afdacf4b6f58bf11c;
mem[1088] = 144'hfb7d043ef824f559f2ffff50fafc06cff505;
mem[1089] = 144'hf478fea8084a07b0053a015809d1f996f4da;
mem[1090] = 144'hf5df09da03c40da20a37f90af6f402d9f0db;
mem[1091] = 144'h014a0e8cfa32f6ac0fdcfdb9f6d510c30c48;
mem[1092] = 144'hf9d7fc810539f3150e5df978060ef0baf126;
mem[1093] = 144'hf30ff591feeb05f6fd8205cfff92f503f700;
mem[1094] = 144'hfc800bd8059a0d1a11740117f3b0f7aefcde;
mem[1095] = 144'h049902cefd53048cfb19f853075ef9280305;
mem[1096] = 144'hfce2fba108e80e6ef4730a5bf4b0fd49fe61;
mem[1097] = 144'hfabdfa67ff37ff39f95cf4f50d29f8c1f485;
mem[1098] = 144'hf89afb600e5df8ef0f27098b08fff22e0631;
mem[1099] = 144'hf977fe27f4fb0caa0164f53df412f6a9f88a;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule