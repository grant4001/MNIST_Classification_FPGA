`timescale 1ns/1ns

module wt_mem1 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h186818cee6e9e4c1f9e4f7b218d90d9f1675;
mem[1] = 144'h15ed1b451144048cf09cf70200270c4a00ec;
mem[2] = 144'h1c61f594e71cff59198a11f4ff39f778f8d3;
mem[3] = 144'h1ea0f081f0c7fc0bfa1e06a3e71206160dad;
mem[4] = 144'h0d2ce356e438ffb10b4900ccfdcee297e5c7;
mem[5] = 144'h1640ebb0e7680885fad70545f7a6fe7fedaa;
mem[6] = 144'hed27f598e06709c0118f067f153f0a8cf86d;
mem[7] = 144'h0c8ded50e4090065e683f9e01edde6a5fc95;
mem[8] = 144'hf9e11248e55c0fb3f449e6f914920217e887;
mem[9] = 144'hffbfe7a2176a0216ff2df105fc351687ed4c;
mem[10] = 144'hfdfb0fb7ebca1a600f1f0640e6a803f9f368;
mem[11] = 144'he874e78509d80e4109020ff2e710f50c055a;
mem[12] = 144'h09f5e6f7e8640e44086fe63201ffe819e91b;
mem[13] = 144'hfda814c50a64ed94eb3318ede64eea7a00fd;
mem[14] = 144'h1cdfee2508c1f059f7daeb7a1a51e550e296;
mem[15] = 144'h1f38f5c5f9f7f62618c6edc51d95fd29e803;
mem[16] = 144'hf4e70343f6e603a6f4970fdd1ea106dbfa59;
mem[17] = 144'hf6e30406e3ff0fb00bb2f2bf13321837e243;
mem[18] = 144'h0f911e83fdacf9c016ddf0bb1d63f88512ae;
mem[19] = 144'h16141e89f51f1d0a02b9fcb40388011600e8;
mem[20] = 144'he9cd1539177ee0d9072de64dfb3c00dc1a27;
mem[21] = 144'he90b1c24f87e0634ee0e01f5190cfe97f121;
mem[22] = 144'h099cf5fcec72e7bce54d0a4cffeee8c3fa9d;
mem[23] = 144'h176e0e5113bf1a25ee2cf96e0c2e03f71e5a;
mem[24] = 144'hf97c0f3c11d3f2cc1e41ec88effbeb001ffb;
mem[25] = 144'h154c170e13e9061c1060196ff69ffc39fc1d;
mem[26] = 144'hf8fcf68a1bbd18b3ed5be6e00389fc8efd71;
mem[27] = 144'h11c0099cf6fb025cedd100f8f128fd5a1e8f;
mem[28] = 144'h1b7e12b710badfaaee241461062a1a8c03f3;
mem[29] = 144'h16721ef30ea5f8ee034afecf07c31b04083d;
mem[30] = 144'hfe30fcfc0f541e2cf570004b1393e40eecaf;
mem[31] = 144'h0bee0fe1e8871a4cf0bae7ef1ac00c4cec1d;
mem[32] = 144'he8e5f3a3fccffef911b5f2a40ab104aa116d;
mem[33] = 144'h016d0d34f3f92079fbf614e9007de3c4f7bc;
mem[34] = 144'hf010f9d40586fb7bebc2f81c0ca216caee5c;
mem[35] = 144'h0c42fe3df1ea080f1cdcfcc8fcbbe57b05c3;
mem[36] = 144'h029c1380134b1b090573e346f33f112bf230;
mem[37] = 144'hfab7f852f4d1f7cce1531ea9ec22fce003b0;
mem[38] = 144'hf6d3ee451809166c057f1a89faaffe771397;
mem[39] = 144'hf1a6f7e7e5f2e47e10b018661452eae116cc;
mem[40] = 144'he0160b6eefa5f7f6f7fa049a1959088f1f38;
mem[41] = 144'hf0d1fe09eccf1812e59201b112dd0383f653;
mem[42] = 144'h18160140fc4d070de34402b2ed0d170e03e8;
mem[43] = 144'h1945f3ebe877feb9e35cf6a2fc601005f8e5;
mem[44] = 144'h159edea80109f5b612ba16daf238000e0ddc;
mem[45] = 144'h0b6be1ddebb0ff9bf59a1334f8beef23f8e5;
mem[46] = 144'h1a3600ee1a9df452fc68e2d1131013550b55;
mem[47] = 144'h0f4d185f0c7b14f7e51b0b80ea410e7ae69a;
mem[48] = 144'h19781f73ffbf0b53e12c052a090ff9bae4ad;
mem[49] = 144'h1d93075b1743f9810d591b16048bf8290fa2;
mem[50] = 144'hf155f28c175200ba0900ed88ef72187ff9ef;
mem[51] = 144'hf3f715bb09edf7d30aedede7123bfa1a07b1;
mem[52] = 144'hea8812a2e3aaf506ed22fabf1e081f87f9a2;
mem[53] = 144'hf7c3111bfe7bfe58f7720e0df5d30c991b54;
mem[54] = 144'h1df3170a0a1bf30019631c110175ec181dff;
mem[55] = 144'h0f7ee59fe24bfc0513000362e36009f90da6;
mem[56] = 144'h15780c1f1db8e8f4e22ce6bf0ed9ff440f5f;
mem[57] = 144'h07a3ea9d1991e3fceec21246f7e5e350f75c;
mem[58] = 144'h077d05ddf5a9fcd705c2fef5e07708a90c16;
mem[59] = 144'he01a0062e00fe9adf81813a901fcf3070827;
mem[60] = 144'he6c018cb0fec02110ad81344ea57162e0865;
mem[61] = 144'h16acfd841e6af0ecf5b106c3006d153feb17;
mem[62] = 144'he6f3edba1c2cf1dfe22ef0fd114afc0604b3;
mem[63] = 144'h0ac9e31812da16b5f3f8f2a2fff309110031;
mem[64] = 144'h1559f64d0fceec750b770125151fe3a41d70;
mem[65] = 144'hfb70f1c7fc920861fa30e68c156703ef10d3;
mem[66] = 144'he90be879f5830e93f1f2fdd10647e12709b5;
mem[67] = 144'h0f8a0acbe957f4f508e8f3871e7e00c8e9d6;
mem[68] = 144'hf878e28fe922e4ffea3404791819fc2618d4;
mem[69] = 144'hebef1925e3e4150311951108f1ab18f01308;
mem[70] = 144'h14fdfdc91ae0e39100df07c4122405df1997;
mem[71] = 144'heb530ac90cdc19d706c8fe41e224f0010ed2;
mem[72] = 144'h07fde4a704cafa3fe6a71e47110c05a91438;
mem[73] = 144'hfff5fd0a1e22f2d0eb9f0d040eebe8171064;
mem[74] = 144'hef321ede026b1ee4f02fe07dfd62048be83c;
mem[75] = 144'h12761047e2f214e5fac1e3e9e1b5fc6d0a4b;
mem[76] = 144'hfb3a1e71f0860828164119a61772e97cf3ac;
mem[77] = 144'hfbd6f5b70e63e599ec1ae83eede11f5f1c01;
mem[78] = 144'h1e810a9ce2bde405174b1151042b1d370889;
mem[79] = 144'h053aec21e3631d44f7611a69f1d81e2ce6fd;
mem[80] = 144'h018d1f8f0000eb8d0416fb8d1724e3181ecf;
mem[81] = 144'hfce317cd1f74e2eae0adf82de941f356f5bd;
mem[82] = 144'he513e4191d0409aaf09af315e256ea62e959;
mem[83] = 144'he6b1feef1b97075cf01d0996fb5416b9019e;
mem[84] = 144'hfca6173201d601a8ed0806f21cd011081034;
mem[85] = 144'h01af06511628184b13bf0aab1c65e3c5e7b6;
mem[86] = 144'h1b5716eeec3be1d2e2b8e0aef9be05c7fe50;
mem[87] = 144'hfba71422f4ad1a14f6b009301c73ed201e4f;
mem[88] = 144'he6fc10f61c980c7bf710189be0da0db0e5fe;
mem[89] = 144'h0524f6b20a6715f7f50cfc2302b81dec14ce;
mem[90] = 144'h0975f53b0f7013ba107bf0751219e13efbaa;
mem[91] = 144'hfddfeaccf0eafb2bf7371fb6fdaa0758ed9c;
mem[92] = 144'h09c10c26f698fc41fae5f36be8b2ea290f86;
mem[93] = 144'h1b64e1dbef580bc1f85201dfe5650b52e811;
mem[94] = 144'h161af3a2077eea38e02b08ff17e31059f767;
mem[95] = 144'hef9200a4e9a218b705f80faff2cffd801a42;
mem[96] = 144'h0c3507030d23f872e11c1e91055bf514fe8f;
mem[97] = 144'hf026ea23e9c1f2c1e9d6f635071717560fc8;
mem[98] = 144'h1813e51310080a890304e886e413fc6a0c6a;
mem[99] = 144'h0156f54ffb0605d6fadff27b1a6efdc9f226;
mem[100] = 144'hf708f5f6e03be2e4e99bf75efee61ffd1355;
mem[101] = 144'hf8a4ffa01db9e371f45b0251e444ecf01500;
mem[102] = 144'h14d9177b06981b551299eeae09161ad2e423;
mem[103] = 144'he6241c2ce0d3ee70ec66062dfd50128612a8;
mem[104] = 144'he118ff00e2aaedc7014b0f75f64fe74901d9;
mem[105] = 144'he80bfa7de9c11e73f04ce1aa036cef930b1d;
mem[106] = 144'hebaafac41f300857efbc19fdfbdeff0e1d00;
mem[107] = 144'h195615b619e30a7e0ace06b30fb4e5d30af3;
mem[108] = 144'heb4bf193f866eca9e2e9faba0f1e06cd1614;
mem[109] = 144'hf27b0d53eccfeb00009b1616fd5e0b751e08;
mem[110] = 144'hf455f56a06b01ad1eb130b1a0b351d4806c1;
mem[111] = 144'h15fe0dbefa76fcc61ef5f6ea0e4febb70641;
mem[112] = 144'h0cd4fe57e7661f390d7cf3dd19730cf0fc61;
mem[113] = 144'h15a107790bd2e875049cf5a000d009730f0f;
mem[114] = 144'hfae80820f55f1c1502a4f2e1f4aa1113080a;
mem[115] = 144'h162bf091e39f0c07eafff0641973f0fc0dcc;
mem[116] = 144'he93fe72ffb3412fc1d4bf5fcfbb5f07afc40;
mem[117] = 144'h162a14b2f34ff011e0991a300330e54d0fe8;
mem[118] = 144'he71500631388f7c00f08e52a06a4e423fa7f;
mem[119] = 144'hf31106b409a7f556ee02e86612a3fdb7fd5e;
mem[120] = 144'hff85eacd0e3ce4f7ea151080ee0a1429eaf4;
mem[121] = 144'h12d5f47ee8520a5a0125f50de8aa0208eda3;
mem[122] = 144'hf41516f6eb860e501f25fbb402d1ecd2fd1d;
mem[123] = 144'hf90bf154f69c13f002c81521110dee851290;
mem[124] = 144'h1af8ec39ff35f054e2a40a6504f3043b1f3a;
mem[125] = 144'hfeee0ed3fdb205d1fb3d15fbe415e1cbff88;
mem[126] = 144'h199ef50b1d61f8f6f330e1fe06aef20bf8bd;
mem[127] = 144'he6c80512e8100f5af12e197fe3eff35f160d;
mem[128] = 144'h0a79ebc70258fca41488ef9df7c3147def9c;
mem[129] = 144'hf3281249198ae01fe703f66fed4a12c8fe77;
mem[130] = 144'hff36fa540880023f1271eaaae64c0b9ae2cd;
mem[131] = 144'h16051e670b3ceaa7189df6fa156a085a0f0e;
mem[132] = 144'h144405fbee5cf4270feb066707ab18b1e4d0;
mem[133] = 144'h0d3c146aef6016a41a820a8fe0f4055d05d1;
mem[134] = 144'heb48005def4ae109e66800ffe1b50e3ef605;
mem[135] = 144'h0e2bfc15ec23e116e3d4efcde6c2e54b112d;
mem[136] = 144'hfa5cf2f808bcef20e7db16010859ff5108df;
mem[137] = 144'hf1041a651a8ffa500473fb560bfd15b71fe3;
mem[138] = 144'h02dffef8e6e4ef88f6bb01f00a31f734e568;
mem[139] = 144'h1d32f26bf4b813dd1a3ff777002017a2e57e;
mem[140] = 144'hf7c300f30e4d12a019f9e80a0241eb6dea0c;
mem[141] = 144'hf5a1e663fd7ef53b1614e3baebf81521ec5f;
mem[142] = 144'h1f24f442f66cec43ff43199716ae0bafeb91;
mem[143] = 144'h0134f63cfd12ec9cea46f86cece21ea5ffeb;
mem[144] = 144'h054ce805014e0e1ff95a1714f61d051710c1;
mem[145] = 144'hfe040901fcd8ee230dc3166de736067a1b86;
mem[146] = 144'hfd7608dffa98f98017a8f44beae20dbb1311;
mem[147] = 144'hf82df0ebf1e809bef5d31394e3120404fcc7;
mem[148] = 144'heba108530a3cef13ed3701a4eebde32fe9df;
mem[149] = 144'h0bd9e90a1bd91cfde63e02c7e8f6fbf8f364;
mem[150] = 144'h12d7ef221731003c128619200588ffe1f36f;
mem[151] = 144'hf88c0f5a014cfaba1222f50c10ace39d1e37;
mem[152] = 144'h1fcff193ecb1ea2f173ef110f5330bbfe961;
mem[153] = 144'h11f21cca1adeeb02ef7cf170f26d0bab17ce;
mem[154] = 144'hf4791f7b03050c731acdef62027bf74f07e4;
mem[155] = 144'hed71e5b116c2e0cc14a7107f19f8f9570163;
mem[156] = 144'h15691a4c1758e5c6ead61ecb061c0d1617c1;
mem[157] = 144'hfd5ee0bffd9afba0eefafe30e998f3590614;
mem[158] = 144'h03c5ef7b0a770fbce3a917fd1c3a17cdf4a3;
mem[159] = 144'hfc61ea5dfb9f1d8e07dee3b8029810c90779;
mem[160] = 144'h1cfd02911d40122ef1cf1f14fa081ef00c6e;
mem[161] = 144'h1a96f5681921fd3114dc1768f0180d8df95b;
mem[162] = 144'h010116d204e50ae91267e708f7c1fd6d1f1e;
mem[163] = 144'hf16a128e11ec1131ed21027df6fe02a2eba6;
mem[164] = 144'h154f12020033f11e0a9bff0a0cd6f53aefd3;
mem[165] = 144'hf3d206b315e5e86c1751e5a916c9e5af056f;
mem[166] = 144'hf8151de319311cbf0d1404c8fae9f737f2b1;
mem[167] = 144'hfc0ef0461b4a143deb26e3831e3f097ff063;
mem[168] = 144'h1fe7f2b30d3e0de5f119f4a4eccb19261af8;
mem[169] = 144'h17750d21e8e0fcf8e9f3ea3a1ae10119139f;
mem[170] = 144'he698071fed2306e11d6e0245e28002651491;
mem[171] = 144'hea4c04c701dce674ea44073f0d96edc9075f;
mem[172] = 144'h175c142c00f8e39b16cbf3320f5eedd7115d;
mem[173] = 144'he0e00cedfd850094033c1aa8eb82e9751172;
mem[174] = 144'he146ee88e149fcfde85df3a2ea2be448ef1b;
mem[175] = 144'h07960b70f24cffccf3fbf119fff0fbb0fd2e;
mem[176] = 144'hf087191aeb7bebf7f4fce112fe2b148d00be;
mem[177] = 144'h1c930055eee8e1d50a1017f1e70818b3e03c;
mem[178] = 144'hf16810de1d68fc321e0b1541e28c1ad5fbf4;
mem[179] = 144'he802ffc71d99f95412e705c3f2f4f925e8a9;
mem[180] = 144'hfa010f230667e91dee0d09f61ec90eb1e512;
mem[181] = 144'he13512d711e5f3411d3be1de092b113704dd;
mem[182] = 144'h1918e97bf0991baaf8cc07dbe2911eea1e4c;
mem[183] = 144'he09ff9ccfdfb15d3ecd60e0ae5e6e7ce1a8f;
mem[184] = 144'hf2f51c7318dc1fe8f4f91d8f16ee0c24105f;
mem[185] = 144'h13eae60fe32019fc16ab12c9e824f9c40003;
mem[186] = 144'h10acf3cd057ee0d11ce7fb83efc8111e098c;
mem[187] = 144'h0c77ef92e4df1735f36716eae836063a0f09;
mem[188] = 144'h18940b841bdbf68aee6202b10b44ef970cf6;
mem[189] = 144'h1474fffe0af2fa6f03a8f1b81398f1ff033b;
mem[190] = 144'h08fcee5ef34e1aa200b2fbfee24600442020;
mem[191] = 144'h17471828f372ebfc135f1dab0409e9d714bb;
mem[192] = 144'he0c6ffc60236f9791198e9a71cbbfa3afae7;
mem[193] = 144'hf9b4f07e15ce17d0f0a4f01c1ff00023fea5;
mem[194] = 144'heed21e79076ae881eb8d1e2f0d641f4bf610;
mem[195] = 144'h0c3ff4870c0cf95ce191eecb0844fae8f175;
mem[196] = 144'hfaf912aaecd0ec68fcc1e273ea77ffeb169a;
mem[197] = 144'hf4b50fe7007ce352175c1d6c151c0ef7ed37;
mem[198] = 144'h0827e7c11363e37019f8e9310a171d1304d0;
mem[199] = 144'heb0b1220178ce561e44d12a7f80bffe6f56a;
mem[200] = 144'h008afa29e4a1f930f20cf5230de8e09a1b75;
mem[201] = 144'hf5d813c7f0780158f17a030b106fe94801d6;
mem[202] = 144'h16f10dce17c41e7f06a30a90091018ece955;
mem[203] = 144'hed4918041fd4e349ea191b5de45a085f04d3;
mem[204] = 144'h040f16790d40e5930026e0d61759f8b4ffbb;
mem[205] = 144'h1c8aef61eebdf31c1d5e13580fddf54feae7;
mem[206] = 144'h14bdffbbf49aece2f3b91a9cffcaeec11028;
mem[207] = 144'h1305f036f3d819380b9ffafae52af5c30c3f;
mem[208] = 144'h0af7f76b15aae2a8e1ccf6551bf4109fe448;
mem[209] = 144'h0968f86fe384e50b1fccfcd3fd1dfccb0acc;
mem[210] = 144'h19921204e9a3fc1c1b8fedf8090b1bafe31f;
mem[211] = 144'h03830768ffde0c4ce28be67ae8b0e8be08a4;
mem[212] = 144'h02210984e8cb15561c2fec28085f02fcea0f;
mem[213] = 144'h0fece0a9053502f90b200ead0cb8e943e38f;
mem[214] = 144'hefc5f38ff5be1a84e7ee0f3511ed0081eeb1;
mem[215] = 144'he5530dbafb011e11125a1e9d00fc0797eb9b;
mem[216] = 144'h15effa9f1c20e1430d6915def500f33e1581;
mem[217] = 144'hedcbf1531c2b16b0025cf3befc5def9eee64;
mem[218] = 144'hf0a6ea5509481a73ef880922eb33e178f6d6;
mem[219] = 144'h1e021be6ea12e091f6d200f3f7f81976e7c5;
mem[220] = 144'h10531039fea400ab13521612e87414baee64;
mem[221] = 144'hee160145ff9eef92ebbbe5871c32f3091303;
mem[222] = 144'h1d240ba0144717170ba205a5081e12d60e58;
mem[223] = 144'hf2f808bcee22edb2e0fbe945e1f9f76d054d;
mem[224] = 144'hfc02f89b0aec005014a0eefdf1ef002e1af2;
mem[225] = 144'h097109b70fa407d41bd7efbc184809fa14ea;
mem[226] = 144'h1a281be115a6030de2e40d30eb24fd8aee6a;
mem[227] = 144'he08be071e657ef3601e90942f7f0f2b31399;
mem[228] = 144'hfb8a1a5de1860fb0053f1b710913ee600777;
mem[229] = 144'hee49ec610589fbf303981901e8f2076aeeb1;
mem[230] = 144'h1464184ce927003dfd76f1f6eb4c0ae61a59;
mem[231] = 144'h09ee0aa918cfe9acedafe659e041ee87fbcc;
mem[232] = 144'h04eefdd107fe0849e19316151c8b030ae0d6;
mem[233] = 144'he6ce0bf5f975f4ca0900194d18d80cba0176;
mem[234] = 144'h0da1ed6f0227feb8ebc5048216c60597fe95;
mem[235] = 144'h08b30cdcf5b9eba0e3cc1135f55c0944f5ac;
mem[236] = 144'he1ee0a4ef74d14ad1902f8dfffbd14da0d39;
mem[237] = 144'hfdcffaca17baf1ede8a6f5200b850129e4e7;
mem[238] = 144'he16617fe02f711a3e5bcf3441fa1f5d7ebca;
mem[239] = 144'hf0220398f060f0b5193905850608e84ef077;
mem[240] = 144'he94c1f42026f0f6c018f0bb213c3fcd9f406;
mem[241] = 144'h1ec1e0f90896e678120e0486f48a0e7defa1;
mem[242] = 144'h06a20f4e0e79f94aef67e27fe3fa19ea052f;
mem[243] = 144'hfaa0e407f26b1cba1bbc1ebb1759e0780abf;
mem[244] = 144'he02806ca1c210f9be974055008bde7df01d2;
mem[245] = 144'h1d22f8a0faeaec98fce3194c0ad013161f4c;
mem[246] = 144'h02f8f1e31212ec4201be17471abde018e26b;
mem[247] = 144'hfbd6f77ff7c711aaee900cbe1ca21d9610ad;
mem[248] = 144'h00e4f406f42deb55e059fc6d05c30792f4b0;
mem[249] = 144'h13681a75f8931740177df771165bfac6ee73;
mem[250] = 144'hfd49ea6fee190702ea310d78fba7e10b03f3;
mem[251] = 144'hee72058eebc0e493108012a303c7ff6602c5;
mem[252] = 144'he514f5220881ee4d0ece01581b2ff9e8e78a;
mem[253] = 144'he3f3f223fc3a147c13eaefb5e5d0127b17c0;
mem[254] = 144'h0954ecccf96ee49907231c07f43ce1f717f7;
mem[255] = 144'he0e0e50701dfec66ff36e4e30d1ced2215dd;
mem[256] = 144'hfe40e3ddec13016416f4ea9df9b7ecee1fbb;
mem[257] = 144'hf2c6e70cee54fbbf05e6f68201eceb3ef249;
mem[258] = 144'hf760f03be6f7f97de0910771fa07f8bc067d;
mem[259] = 144'hfc1a1ae0026fe8b0068be682f0041bb1f252;
mem[260] = 144'h0a8a0f220c83f105084ae0fc1f2fff0eec3d;
mem[261] = 144'he0fffc15154ded19f51d12c7fddb147f1396;
mem[262] = 144'hecd4064b1851079807171316f4bfff4b0379;
mem[263] = 144'h091eeb79e87a00280eabe8b0fce10ffe1aa6;
mem[264] = 144'he1a3171b03eb05a8e5361b7bfb980228f297;
mem[265] = 144'h00c4e60010d301601e34f500098fe9bdf4a0;
mem[266] = 144'h0102f478f33af34e0fb5eb3d1ce1e2faeba6;
mem[267] = 144'hf08805671d4b0d531fc10781e6fbe745f812;
mem[268] = 144'h04e4fe55085606471a4ee78ced46fe40f169;
mem[269] = 144'h12b5094d03be1af0f40af182e689f5720247;
mem[270] = 144'hfd6cf8d6f080ee97130819dffe3518390e50;
mem[271] = 144'hf22c0549f94d0eacead9efd901a80178f62d;
mem[272] = 144'h1437fdade86f0d100ca7efc31ae4e1e6086f;
mem[273] = 144'h16a6f34a1e2f01c0f2cce1bc0df01fe80523;
mem[274] = 144'h064f0e08ea5410160afb0ad7fda20697f029;
mem[275] = 144'h122f19f7e0b700bd0679ebf7e1bd06efe90c;
mem[276] = 144'hf06f0da60379e742ebcbf2ccf8c317f010a0;
mem[277] = 144'h137e1902e9e6e5c5e5ae02061b27f811e27a;
mem[278] = 144'h16cdf0f8150c1802e31ffe5ff19e01f20aa5;
mem[279] = 144'h00e2fbf7fb7a0e690dacf46d1f18f8d6002f;
mem[280] = 144'he083035fe57c01ebf289ea43ed18e164e758;
mem[281] = 144'hfc46f2f9ea2c1a8904a007031e34146eed87;
mem[282] = 144'hf4ea07f4f78110cdfa4de3170731f83f118e;
mem[283] = 144'he3dc030b1accebf20ca00c381d4fe8530c3f;
mem[284] = 144'hf6c9e3781964e569ee5114b11413fda9fd75;
mem[285] = 144'hfecae2ade1861182ecaa001011780587e403;
mem[286] = 144'h06f6030c05d8e1bdfdb10247156e0f7af906;
mem[287] = 144'hf8cf0423149e09f20c75e16f1bf40e02f479;
mem[288] = 144'hed58ee68e7ad0eb2f8e308100493f478f4b7;
mem[289] = 144'hede6f2ce0d85155e070ae2e2ead5e895e3c3;
mem[290] = 144'h0ac90c63f302016e19e8e262ecf903dc09e1;
mem[291] = 144'h151f1538f21ae2a70935e09a1ff71914efb8;
mem[292] = 144'h05e20c29f2e8e322e54ee2e6f0c0090d075c;
mem[293] = 144'hec971b8ce6fee04af538f5da18a513d602b5;
mem[294] = 144'hee161a82f883fadfe1581e310d0af38b1b91;
mem[295] = 144'he86c1412f8f61205eea8fa6deee8f2cff7fb;
mem[296] = 144'h0b080362efc7f5fa1705e095ec0f0247166b;
mem[297] = 144'h0561114b164cf1d710faec7c174ae626fe98;
mem[298] = 144'hf96de3fd1508f544ee471f9508340b6a0474;
mem[299] = 144'he378fccb1bdc1362f414f690e684e53d1cfc;
mem[300] = 144'hf43cefef0e1de295f97c1760fdd9e792e650;
mem[301] = 144'h1930f613042a1cb0193ff93ce01b0410edbf;
mem[302] = 144'he558efa9e06a1f1113e1fcd1fa44f948f4d3;
mem[303] = 144'h184d1aa71eb6136c086ae0ca1e56fe0eefad;
mem[304] = 144'he0960a8c08d01de2e40808a31cf4ee02ea4a;
mem[305] = 144'hfe320c9fe500e4fee5d5e1f7e9e80b1d193b;
mem[306] = 144'h1941117efb1cff6304a2e03717a71623e3d9;
mem[307] = 144'h05c51a7a05b2f3ff1b0115b206f8fb000c49;
mem[308] = 144'hf6e71adfe2baf1acedb112ddfd4dfcb0e9bb;
mem[309] = 144'hf07806d1013eebfa160ef1db0d4fe37ef0ce;
mem[310] = 144'h06810618ec3b1b8ee70201bd1cf616031ed8;
mem[311] = 144'hfb8ce9de1f141cf2f95ae15ff7211966115b;
mem[312] = 144'h1683e54af6410dcae5aa1587e05de0e61e8d;
mem[313] = 144'hf42b0154f5551b440d3df502fe6b1774fff3;
mem[314] = 144'h0113ed1e14d7ef920c5517d9172b014e1fa9;
mem[315] = 144'he084fc9ff9ea00c3f5dfe4c5f8071a771f84;
mem[316] = 144'hef2a0f7df56c1c6ce91e15a5ee900eddf4bc;
mem[317] = 144'h13111e73f482ea5d1cc9e6fe14c4edc80a59;
mem[318] = 144'heed506d016e10bfcee3a1d06feaf1e6af6b8;
mem[319] = 144'h13d3e83cf4c6fcde17a00f2319231cb2f656;
mem[320] = 144'hf34a1624ea99107f0f8aec37ec691b2d13a7;
mem[321] = 144'hf280e2ea0e0b04c2f0be10b2002a1b9808c2;
mem[322] = 144'he5970fd201d2e5ade9f3e91e0644f23a1c31;
mem[323] = 144'he9130b6feafff498ee08feb6ef90f98be490;
mem[324] = 144'h03131e0d16a40a1201b10d87e752e8c7fd19;
mem[325] = 144'hfcb40e9f035909b0e53afe58092be5bd007f;
mem[326] = 144'hef78ea5400ba01ee0345ed4d1495e3b6eae6;
mem[327] = 144'h1f94e1521eb106f3059507a0f0e5f8b7ec25;
mem[328] = 144'h16bdf689174ef66b1a36f5e9162014a001f2;
mem[329] = 144'hed010779087a171a1ddaeb551a0300e91549;
mem[330] = 144'h024d09a704b3f87dfcb40ff61aa91bc31f73;
mem[331] = 144'hea4c0e75f0280fc715000888e0460c5c108e;
mem[332] = 144'hefb8e54d160ffd1ffdd6077fe61501e7febe;
mem[333] = 144'he91be53dfeb51b25014119e6f57711a5ee48;
mem[334] = 144'hf462f1630401e9dd0e11e7abf9cb11f8eadb;
mem[335] = 144'h1f1ffbb6f18901a01c2f04f20196e641eb2f;
mem[336] = 144'h13120414097503b61a3110b2f2d812321875;
mem[337] = 144'he932fde7fa70f0a6fcdae267e462fb31fdbf;
mem[338] = 144'h027ff460f19bf00e00271732e1790a74e5ec;
mem[339] = 144'h05f811bbeae31cb118a2fdfcfc0b0373ffea;
mem[340] = 144'h11f7f50d0630081c0aab0254f6ebe9090ba7;
mem[341] = 144'h054a193dea7a0620e8f4e08df06b138e0541;
mem[342] = 144'h19bc1ae2f1c8160b06b9ec8ffd0a0231e031;
mem[343] = 144'hf85d13c1f3adf37affb0000ee0d9e0c6fe87;
mem[344] = 144'h1071f55de65c02c3e93ee80bf1f210140352;
mem[345] = 144'h08d0e7a0e200f4160839fd55f4d1ea7af625;
mem[346] = 144'h1e46ef20e098e3c6093a143603531d371c1a;
mem[347] = 144'h0575ea10186d032eecad14fbecf90297037f;
mem[348] = 144'he9a403cf00e91d0cf8f5f45504430eddf063;
mem[349] = 144'hf520f7c91d53fab30094fa6a17dff9e9097d;
mem[350] = 144'h111af88cfe760c5bf71d042718a9f1f80fe1;
mem[351] = 144'h1a4301c407ab0fc3eb1301f4fec418131227;
mem[352] = 144'hee5c10a8e48a09611cb5065d1144f84d05c3;
mem[353] = 144'h0d1efce71c7418aaf069031719f1f9f40082;
mem[354] = 144'hfb6c00ab14fdfca50456f1ab1990068bf560;
mem[355] = 144'h0e7a0c650b49ed45e3201a260f0c06291f1b;
mem[356] = 144'h03c5e611e13004befd60058e12431ee3f200;
mem[357] = 144'h05f6f73ae98b1c4ef263fb2c0d180310e2ea;
mem[358] = 144'h0902e6dae68e10ac1223e13ffa8de091e7d4;
mem[359] = 144'h15bbf6991bb019551d43f618e488e8900535;
mem[360] = 144'heec915d10f40fdff0b2f03caf9bafe230257;
mem[361] = 144'hff1e03ef0858e8010303134508d60fc6e2d4;
mem[362] = 144'h1f75eabffba205e4145115f414761436e74a;
mem[363] = 144'he588ed01ee36e08ff181fc40156f0684e5f3;
mem[364] = 144'he7fb1d3d126513dc11f01fedfee4f109ebda;
mem[365] = 144'he48c17ade57cf50e195e1bc3e0d3eb2ee772;
mem[366] = 144'hf600faa2f4260b7101c6ebc319c4e1ea1178;
mem[367] = 144'hf70b0bffe62eeaa8f6fef90bee2fec59e512;
mem[368] = 144'h15140bbf1c9ff3e5e8dae37ceb49efeeec22;
mem[369] = 144'hfef2010cea6aec28ee7d1fc9051fee2dfc54;
mem[370] = 144'h077f117a12bd08d4ec0d0207fcfd0a0309ab;
mem[371] = 144'hfb6becba0474ff5113f8fab203b6006719ea;
mem[372] = 144'hf34f139e1bb9ecd3edcaed80f3871e3307fe;
mem[373] = 144'h1ddced08e3cd08f914fe0df70f0919431803;
mem[374] = 144'he96ae91febfe09881d06f5fd1f6c0a76ea6d;
mem[375] = 144'he31dee27132bf6e51921e0a0f849087816dd;
mem[376] = 144'h0181f36ef20fe0d5edafedbf0e08114ff4de;
mem[377] = 144'he6911d3611cc0ad403f9fbe21bdffb831379;
mem[378] = 144'h1376f0b60995f155196318abfd3ffa76fb36;
mem[379] = 144'he427e161fc74f32af8bfe4f60be1ed5b1cad;
mem[380] = 144'h040c1c63fa16fdf0e640050f0cabf1ca0899;
mem[381] = 144'he510fea01c000489fcdef7cfefbef399e71e;
mem[382] = 144'hfea8ee04e30d1e3d05e6e614edb71aa5fea8;
mem[383] = 144'h116807490d16e8d2e3d2e93ff5e9f2e3f820;
mem[384] = 144'hef1c04c2fa53fd1c1b9de49be132f3e9ef39;
mem[385] = 144'hf0e7fa30fb75e392e0dafb6a0edf1ccae84e;
mem[386] = 144'h03c504a9f1850d68f4c0016ce3b7f3d60040;
mem[387] = 144'hed94fcff0350fc76e21602d8fc3105ae04d3;
mem[388] = 144'hfd7b0bb2e0a0fa33ee19fa7e0ec3fb731c45;
mem[389] = 144'hfe630209fb65fcbf0386fa6110d4ec07fed3;
mem[390] = 144'hef61086fe7c51b7fec78154af2c2028c0418;
mem[391] = 144'heb6f13ed1c0ce79c0e750c660421033d0af8;
mem[392] = 144'h00c6f558e7b5e86df4ca0a3716cd04f60352;
mem[393] = 144'he4180e9bfc1f1230ed04e577f9e8ea1d0b96;
mem[394] = 144'hef17f0d4e359e92418b70bd31e23e527ed8d;
mem[395] = 144'h028c18b0f7b9e7fd0676e5da0e17197d0a7e;
mem[396] = 144'h01b1f7941734151cecfc0cc0e15b090c1f32;
mem[397] = 144'h168fe58b121ae160f891f6711280132c17f4;
mem[398] = 144'h184fff6611601387f1fbe76901ce0872151b;
mem[399] = 144'h1a130ba5e328186efd50ff3309ab11831587;
mem[400] = 144'h0faff2b707d7ed61e1921e131a82199002a3;
mem[401] = 144'h0b0e0e23e2ad008eed0df1f9f56d059711f5;
mem[402] = 144'hee741d0c07671f870dd30454e6cdf53901fa;
mem[403] = 144'hf0f812661ddf1489fa900cb806a2e87210fb;
mem[404] = 144'h1af0eb160905f23218f70103094910630447;
mem[405] = 144'h07f51b97ff41f81ef4730632f9741536ec1c;
mem[406] = 144'h11edf058ef5c0ca8fd77f12df391fb5b039b;
mem[407] = 144'h0d25e6e007c2f71de5c8f62ceea2f029ec86;
mem[408] = 144'h07df1334156c0c870033fa60fbcff438eb67;
mem[409] = 144'h0e411b46e6e6f8ae0b1d04f318cce549149d;
mem[410] = 144'h1c730fbd0db5099cf4bbf9d9e05fe02b1903;
mem[411] = 144'h14acf099f89707ccf1a5e6ba00a503bc15b2;
mem[412] = 144'h0fffea460be3ee0713b41f350dc017371534;
mem[413] = 144'hf3e51eaef9affbfa036d0799ec9519b8f45a;
mem[414] = 144'h08a3ffcee222e4a31c1c1b000cfcfb7c03e8;
mem[415] = 144'hf2e514dc05fe097ce5cb0fc6ee51e3b418be;
mem[416] = 144'he253ed06eb6fefede11df487dffa16bc18fd;
mem[417] = 144'he4710de7147bf4850322f942f97ae9f5ec56;
mem[418] = 144'he6b0eafbe6801ba90363f5501fe6ec0bf844;
mem[419] = 144'h1f90e0200838e11e060fe50feb9510be0fcb;
mem[420] = 144'h18b7fec9127a1562f34d15a715b803c00c5c;
mem[421] = 144'h0780ed70e056e09011e605d1e3fce4021ece;
mem[422] = 144'h17bee0a3040cee9d1a500a16fbc5122f107e;
mem[423] = 144'hf310f035f78afbf2f4331eda05d1f9671bbf;
mem[424] = 144'h004e066f10e9f993e040fab40da7f7510227;
mem[425] = 144'hef83e36ae557f8c6ebc10375077d174be87c;
mem[426] = 144'he258e7f904b71ad8ecfd1d7ae5f902b1025a;
mem[427] = 144'hf6b0ec40ec4806ace02efda304a100a51e48;
mem[428] = 144'hea4be5c6ff871c31e02803cf04d0feeb0672;
mem[429] = 144'hec22f645e310f779edf7f0370cb2171f1ed7;
mem[430] = 144'he42af04dff491ea9faf1e58714c7e2031b66;
mem[431] = 144'h12f500830e191f64113514bc0611e4c4fe7a;
mem[432] = 144'hed87f29806711d87f8620575fcd9f9d606f1;
mem[433] = 144'h0ad5e83ff58e186419d116870779e7eb13df;
mem[434] = 144'he0a31a100ae1e5e7e91bfa751772e6721136;
mem[435] = 144'hfec2038df4c51277ec98009a13bf09aa0c80;
mem[436] = 144'h18491c1e01b21078f0010a3c0152106d1ea1;
mem[437] = 144'h07831ed2f0bbedde18281ea10ccc065a19c5;
mem[438] = 144'h031b167a0e9b0d05fa9eeac0fbc4ea1be712;
mem[439] = 144'hfb161389fa320d38eb901441192feb290655;
mem[440] = 144'hf409e6461101ee22e2e50d6d18c4eaaaef12;
mem[441] = 144'h0cdf0e6507fd1682091ce24ae5bf11b6e38b;
mem[442] = 144'hfb2bfd36e6461b27e379130319360723e6a5;
mem[443] = 144'h014915a4f0970bb9134a1531f41de721eb19;
mem[444] = 144'he90a13f60ee9f2f3197afa440430eba7ed06;
mem[445] = 144'h092ff961eb2f1a5ae13dfabbe56d1b481e67;
mem[446] = 144'h050efbfafea404ecee6a0812e992e689f906;
mem[447] = 144'hff59e98e1984f519e275fea5fd03f450ffce;
mem[448] = 144'hf18dfb1205391aa40d6f11cafab906e4eafa;
mem[449] = 144'heee107d3e2201afc0bc312c1fa7b12141abd;
mem[450] = 144'he3c91024f63c1d07f858fa85075ff257f215;
mem[451] = 144'h14f9fbba0158029c12f3ff29146bf6780b59;
mem[452] = 144'h1e1ae8d6f2a4176b1962feccf8691e75198b;
mem[453] = 144'hf7e4faa5f5ebfc5d0488f1a9f94ee3d7082c;
mem[454] = 144'h1906f3ad1065ef3cf312f282fe37e9b30eff;
mem[455] = 144'h0228f37f0e0e193fe6b3fbf009a910ce09d9;
mem[456] = 144'he1f20fb4e611e72a18811ad30861f76afce3;
mem[457] = 144'h02f9e543f418fcbefc03ea8b0e0df11415ba;
mem[458] = 144'hf94305c5041bf4de16be0b951768172cf02c;
mem[459] = 144'h0205e8961d12e3fbe07aeebcfae91bd31ae0;
mem[460] = 144'he6d10b97e5b71ae40479e0da1f9d0fd5f114;
mem[461] = 144'h0d4a07ea1aacf183f7b5f5de14db1367f9b2;
mem[462] = 144'hfcc1e8a50072fe5aedc5fbad0000151df74d;
mem[463] = 144'he5ae19d9ed0f0fb6ee16e1430dadf03a072b;
mem[464] = 144'hea1fe8fce1f7e5490a231461ec2dfe95fc68;
mem[465] = 144'hede7e694fab5f91af6c2161a0b0af380f052;
mem[466] = 144'hf4a7f2510ad9ea6bf9611ef9e1baf6b6098e;
mem[467] = 144'h06a3e3c1175ce2e9ed8116c9ff37f40bf214;
mem[468] = 144'h10260a380837faafe7aa169407a2e2ae0981;
mem[469] = 144'h0c39f130e0c7f5b803d0e2bd1565eee5f797;
mem[470] = 144'h1c5a19d1e9410296f060f714ec2c13cb0203;
mem[471] = 144'h114c0cdd0888e707f1ea04ad004212c1f805;
mem[472] = 144'he2b7f6160d79fba2e45f09181f1a1716ef8d;
mem[473] = 144'h110b0e4f165215070afc1ae9e80ef21d1283;
mem[474] = 144'h05fc15ebe9dd1b9814901b54f9f0f6cb18f7;
mem[475] = 144'h169b0b75f7851b39ecd20d681ce1e5961576;
mem[476] = 144'h1be7fd13e8ddf3b3e98c1f00ec1e02bb0369;
mem[477] = 144'hfb8701060874f7eee365fec5fbaefa711da7;
mem[478] = 144'h1f460ae00132ed39f76ae2a50180fd7fe6a4;
mem[479] = 144'hfc031d5708ea1d40fbfcef250dbae281f7a0;
mem[480] = 144'h0e2900251eb9e58d036bf1c6ef1a1654153b;
mem[481] = 144'h1d9814d5f1cdf1b7f0e2ebb31a520e201bac;
mem[482] = 144'h11e30827f2e61e1c04e9e3b2f4a4024a1b05;
mem[483] = 144'h1456fc411f9c00e3eb290750103bf1860540;
mem[484] = 144'he0ffec6bfb3b0f850a92fed106b4f6771ee8;
mem[485] = 144'hf35f0e870cf2e8f80daf183cefa1ee3c1b8e;
mem[486] = 144'hf323fd55e7e1f829159f0a5fff761f68fe47;
mem[487] = 144'heee10b19049617d41fa81e6909a1fea7f501;
mem[488] = 144'hffadf111fd98f334064af56beb89e30a16ca;
mem[489] = 144'h0e9fe2d6e533157b15eaf8dc168207021f58;
mem[490] = 144'h1c401774fd18fae8e73dfb5df4b01634f08a;
mem[491] = 144'h14011de2e026092a023c084f1bf1eba6f24a;
mem[492] = 144'he0b204c00c5510450e7c049bf85cfc57e27b;
mem[493] = 144'h17cbf941f7f51a70133b0349f426f429e730;
mem[494] = 144'he8950286f36815f5100f1e85fbd40cb7e7e5;
mem[495] = 144'h044e00d0e2d91177e9c41b64e45e13690f61;
mem[496] = 144'h013702be054c090c11050d3a065812201573;
mem[497] = 144'h1a3417ac1d78f24e16bc00f618d7e792f90b;
mem[498] = 144'hf578fd9f0b8c0635e13ef961fdaf1f6af52a;
mem[499] = 144'h1d2715bb15a9fc850749e784f9e1e992079c;
mem[500] = 144'h1f83081802f8e47af4f5f16d0247fe81ea7c;
mem[501] = 144'hf83e022e1659e5a9f54218d51d7bf0921982;
mem[502] = 144'hffccf509ea9d08810c75044f17d7f25b060c;
mem[503] = 144'h080af2021420e597fc1b1bd9109ae57be20e;
mem[504] = 144'he36eef40e60708e9f5cf0e0908361d8ce33d;
mem[505] = 144'h03e30577109d1920129e0131e338e305e1d1;
mem[506] = 144'h03360de50e7805b21db0ff94eeebfcee165d;
mem[507] = 144'he439e1ba1eab12bbed3d0e7c018a06ea0070;
mem[508] = 144'hed0b1a320e06f6290df8f41b08bfe5831e13;
mem[509] = 144'h194e1e0af462e49f1384f3c1159ff5f9f47f;
mem[510] = 144'h0bde04ebfd5c06ba1cf4095406d2141af079;
mem[511] = 144'h04800bb01f950961f201f1d7fd7ce7ac1c3b;
mem[512] = 144'h1b66f4a3082a13a4ec90030f058af8590be2;
mem[513] = 144'h1eec1c26ff39ea74e867fe6be8a7e86ef5ec;
mem[514] = 144'h07a7e848f934ef6004f712a5e656e1ce140f;
mem[515] = 144'h098f0786f634ff721c3a06d40e6ef5581416;
mem[516] = 144'hfd2b07baec361d57f4df0ecc0ebaeb3200a0;
mem[517] = 144'h1099f7f4fadde03d1bebf7f719f205eae34e;
mem[518] = 144'hf89c1f5cfbdd1f2ee05a0144eb63097d1ed4;
mem[519] = 144'h0deeec9fe960edc9ecd90213f4e2078bfbf7;
mem[520] = 144'h178216320563e53f1a75ed6e0ba7e0e6ec37;
mem[521] = 144'hf159f32c0c49100510d4f470f70f1531105a;
mem[522] = 144'hf09f1632f60dee091351fcecef421064eed7;
mem[523] = 144'hee8e028fe75f036b1da4edde0f69e5b40b43;
mem[524] = 144'h091419da1767edeae4780f03e81305caed6c;
mem[525] = 144'he95ef098e08ee6a3034e1ee1fc91ff431fc4;
mem[526] = 144'h14a0ef5bfc5bf52b01a706b801bdf2dff451;
mem[527] = 144'h1e88179ee329ff82ffed0ca9f67014b3187b;
mem[528] = 144'h00581b11f151198dfed3ec37f7e0f50416e5;
mem[529] = 144'h164fe773e31602dff48613290f791f73f760;
mem[530] = 144'h1f8b0329f914e4801ba90607048b0d691269;
mem[531] = 144'h082a0f740ff50a3c0a57ea81e9d8154de105;
mem[532] = 144'h0150fc390fa60bfb14d51e0cf816f6c70826;
mem[533] = 144'h007bf87f1404130de784e9cdf47f0ca3e5cb;
mem[534] = 144'h1cf814a3f32f11b908f2e452e08b144df7bc;
mem[535] = 144'hee01f13ff10ce07b0f961aee03781e5d1490;
mem[536] = 144'hf56d042d1487e5440a89f468eb00ff52193c;
mem[537] = 144'hf646fa990d170b2d031a024517e71e22ea97;
mem[538] = 144'h09d8e8ddf30a1edce50ce0b71d36152a0e2a;
mem[539] = 144'hfc880941f337f84b0062f5d9fae7ec57efcf;
mem[540] = 144'hfb11e7eaf4bce02901d5ec790f980b4ffe07;
mem[541] = 144'hf545ec0e140f0a8eff6b0378e58016670a5d;
mem[542] = 144'hf867ff050b660cf9ee090e36e365f3fdfc2a;
mem[543] = 144'heb33f061064e152307effadcfe4c0c0ef59b;
mem[544] = 144'h16eeef54f4b2fbf4ea76ed9403f31409080e;
mem[545] = 144'h03c9f55b017f0ec9ee5706fef04aeadbf7df;
mem[546] = 144'h09791e0ced3ff334e6d7f3d0f4db19eee7f5;
mem[547] = 144'h09611be21c1f0058edc1f98a0095eef3edb8;
mem[548] = 144'he5b00a2ced9ff0a40337f80ae7cb18dd1333;
mem[549] = 144'h075dede61f5bf2cb12d3eabf111b1b04ef45;
mem[550] = 144'h1c07f2c402ba0de11400115bedb0142ef1a0;
mem[551] = 144'hff50ea33f7f8f9441e6f10ad10b4001109bf;
mem[552] = 144'hfb16eeeee950135bf175ea78e971f87111af;
mem[553] = 144'h10e41d5aea60e7b3e0b40b9a00fa1001f3a6;
mem[554] = 144'h02bde897e2701ebb0ce91c4907aaff13e9d4;
mem[555] = 144'he91e0f76e2e41655e35f07c81c67e3870d2a;
mem[556] = 144'h1d4ce5dcfff41ffbebf5f286123211380d67;
mem[557] = 144'h00c8e7a8009a0a3d0bae0763e6c8e691fa39;
mem[558] = 144'h0715e9eff3e10823f5bf1d2f04d10501ef52;
mem[559] = 144'heb8e100cf2f905c7119ff2021d83f955fa11;
mem[560] = 144'h0c01f36ffe73114419e2ec2be406f8c6f774;
mem[561] = 144'h1e98e4bc197a0f23ee231655f79e0d2c0142;
mem[562] = 144'h028cfc4c0e5f14110edc19b7fcd5176aea13;
mem[563] = 144'he3faf4d20ac20f7b1a7802120ac1e46e1f3a;
mem[564] = 144'h123ffc9ee6680f150944ef45f77ce46dfabd;
mem[565] = 144'hf9bc1617fbba0d87f51eea6d105909f5f567;
mem[566] = 144'h0ef718131b2d15ee0a56e1f002c0f38af502;
mem[567] = 144'h18b3f0b1e6990b2300481ea3e9b2fe741fa5;
mem[568] = 144'he032f177177c0f62f931ec51e91f0bf2e897;
mem[569] = 144'h03deecb4f4f9e1e413ccf53405921b27f74b;
mem[570] = 144'h10b4f0dc02a8ef8713351218e3a90421e4a8;
mem[571] = 144'hfc0f05b104cd1dff1c7bfc160d5616a4e838;
mem[572] = 144'hf22af19c0a99fa9fecbef4dbe0b714baf9ae;
mem[573] = 144'h193808320a6a14f01daae1491edc0411ed88;
mem[574] = 144'he0bde7abec1fef79f21a1750e4890e1916c9;
mem[575] = 144'hea041defe0aef1ceec74f17c0f7b0771ebd6;
mem[576] = 144'hee0c11de1140031bf1b6fae4e13e1282f22e;
mem[577] = 144'h19abfcbd1f3414071684120d020307730cea;
mem[578] = 144'heedd05d21470e4e91e1de5f604fbe7a0fa8f;
mem[579] = 144'h1c0c0fbefecc1c68f8551804e9c4ffaa1450;
mem[580] = 144'h0def1681195efea21617ef8813e4e5f0e382;
mem[581] = 144'hecace4961d94fc62e7550618062d086d16ac;
mem[582] = 144'hf652f3f4f02bf0c3f56a0b5501a1e44218d2;
mem[583] = 144'h1ff9e7650f5212881d4cfac01a7e1ff30665;
mem[584] = 144'hfa3c190b1e0ff8b6ea0716b0e5cf039ef6d8;
mem[585] = 144'he75eff9410220745141ced250cd9e6c3fb48;
mem[586] = 144'h0b94f075edfb10bef40a1d8a0d18efa704ed;
mem[587] = 144'h1c7b19d8f700e4fef38cfee4023e13d1e4d2;
mem[588] = 144'h18ca013ee59209ab0c5e0c0213bf0019f075;
mem[589] = 144'he01d1da91ef9e9dc0b671a6f071bf02e1d05;
mem[590] = 144'hf2e01253eb000646e07ef6c20307e279f348;
mem[591] = 144'hf3800c5112821321174c1bdee4d30ef8fb6a;
mem[592] = 144'h0cb4e7d1162d0e2ee414fa5be1e5038119c9;
mem[593] = 144'he6ee096feb30eba8e702ed0f0a19082ef27a;
mem[594] = 144'h0f5ae71b1b4bf6b006f8f46be4cb1d240bfe;
mem[595] = 144'h198c17eef2591328e23e0a35e410e7e4087c;
mem[596] = 144'h02e80d4514a117c50615e1371974ed2c013a;
mem[597] = 144'h0075f787fbe3f2f3030b1691e977f9cce11a;
mem[598] = 144'hf6d01e18066bfd8b1d7018c711e907b611fd;
mem[599] = 144'h126d0302f4df01391aeaebc30f180e04012b;
mem[600] = 144'h0c9d00f2e6201f200fafeb5f1ab8190e02fd;
mem[601] = 144'h064ee5ebe76a0ece09970aa917a21a151a8a;
mem[602] = 144'h00dfe8951e1fe29408130119f1001b2ff614;
mem[603] = 144'hf3421b5c080b0adeff5cf0891fe011b1027c;
mem[604] = 144'he432f67811570eeef44210ff1cc9f438f103;
mem[605] = 144'h1d7503c41aff0dcb092c081cf273e83f0188;
mem[606] = 144'h114ff9a0e07e19a5f976f6b20385ef2bedae;
mem[607] = 144'hf4ae126cf916eab1e122f436011e0da6f4fd;
mem[608] = 144'h01a3041a1b5ef7650764f424e58602c40e4f;
mem[609] = 144'h00fce1bbfe82f7860e42efe9f6dee148176d;
mem[610] = 144'h18e5ecca00e7e8730e0f18c4e3abfc380a18;
mem[611] = 144'h0c76fbb90615fc04ee8d1268f591f9c20ba7;
mem[612] = 144'h0fa0fb6d1880f4a4f52f1ee4f631075fe89c;
mem[613] = 144'hfdade6cbed42f0c609a5e2c4e2aef705f08d;
mem[614] = 144'h11b61b16ef2ef739024cf7f90882e943ee9b;
mem[615] = 144'hea3e0a2c0619038e00eb18b91a0efdb7e49d;
mem[616] = 144'hfb1e1366f8cf06b8e24ced9516a0044fe8b1;
mem[617] = 144'hfa45159617841cf5e3701c3fed3914b510d2;
mem[618] = 144'hfb6c1744e30804ebe77116d5e8bbfde91bdb;
mem[619] = 144'he635080c0cdbfba704171b51edf7fde60b65;
mem[620] = 144'h15fa079b13c00f6c1754089cfda50f53f420;
mem[621] = 144'hf3e9f389ed11e737fb10fae9e3b6e6a51bfe;
mem[622] = 144'h0a55ffd81d9c0ecf1a5e043f187f00a21857;
mem[623] = 144'h15c90cfbe22bf85be37be616f21eebc104db;
mem[624] = 144'h0d8f18d70fdf1ddef77afb0106fa01f2ed26;
mem[625] = 144'h04501036099319b01f0e10b901ce18fa14c9;
mem[626] = 144'h1707ea6eec5cea20f3600a14f343180d0b85;
mem[627] = 144'hf3e60174f58ee5c81a0be813fc93e5e213c2;
mem[628] = 144'h0bfd07b1e5a403e8ed88135ee105f180f77d;
mem[629] = 144'he8a81a76ecebf19e0743059a1703fd220e36;
mem[630] = 144'h130fffe6f5790781043706f50b93141e0985;
mem[631] = 144'h0841fc401916ff98f69c1e9a072ce12e0a68;
mem[632] = 144'hee4d19dd1143f72f1e8a1044f7160d4103f4;
mem[633] = 144'hfb3809350365081dfc6be86ef89d09540a63;
mem[634] = 144'h1617054000ff0cdbe54a0936097d094ce2a0;
mem[635] = 144'he2951a1718c807c619a61161f5610c6b0c8f;
mem[636] = 144'hf1b617edfec7f19304c1e68a0ee0e6341de2;
mem[637] = 144'hf69f194ef58217d60a25e562f9910c9dfc62;
mem[638] = 144'h1f6ff4b9e7d7089cebb2161ee31aef96fc1a;
mem[639] = 144'hf0dc1a61e7a5e04fe677e6cbfad1e6610e03;
mem[640] = 144'hec0e171216c4fefe160f1154eeecf93fecfc;
mem[641] = 144'h09f4f365e9b91abbfb0e12d0f3b2e54ff71f;
mem[642] = 144'h0636e25c0696e3fafd610bcf0163175be09a;
mem[643] = 144'hf5f509c01d671bc0179d0194105a0e12f1e2;
mem[644] = 144'h071f09090cd0efbc080b0410e1d80fdc0c95;
mem[645] = 144'hfdb0e267106fe4b71025efd205a815ede5a8;
mem[646] = 144'hf600ff9c0a92f3cce7790c0b0c851ef6e206;
mem[647] = 144'hf4d9ff34f26a1bdd08b916ba083f00fcfa3f;
mem[648] = 144'h17fd0ca1f2dd10b2004e1652e5f60079fafd;
mem[649] = 144'he7c3e06417cafe01f320f38912fc2033160c;
mem[650] = 144'h0f7b1c39e03901eeed6eea32fdd01b7118e6;
mem[651] = 144'h042f0ca7eaaa05840cd8f43405aaf048e5c7;
mem[652] = 144'h0491e0b2f6ede971ecae0abff357ed370561;
mem[653] = 144'h0411f43ff50503ec1ac7f1caeb571847e566;
mem[654] = 144'hff2df838f420ed150187ea6e015cfb1e0521;
mem[655] = 144'h1bd4efc8e3f1fcfb0eadf4691995139519ca;
mem[656] = 144'h04a5ec1000efe9f610f714fc1199135ae925;
mem[657] = 144'hf617fa6dffba0eb209721c2e08c0188909b5;
mem[658] = 144'h09e8f174ecaf0cebe313fe5503f6f6bbe83b;
mem[659] = 144'he4e2fe00fc49f83705471990e85bf5e80a85;
mem[660] = 144'he54518d1eae5e89cf0d6f8e31661f391e84b;
mem[661] = 144'hfeb4ee8e1c3e12b3ea67eda6e527f90116f5;
mem[662] = 144'hf56d1ee7e3590879003211d9ff24192c1de6;
mem[663] = 144'h064c1cef0f751912f181e307f6930c6cf0a2;
mem[664] = 144'h1653ff63180b0dfb0a81f494f5120943f813;
mem[665] = 144'hf5b81d371e52ff1cfba90f62ffd1edb6e3de;
mem[666] = 144'h019effd7115eff58e9d90410ef83f644f540;
mem[667] = 144'h1dd2e141e109e9320700ffcf11a30cbaf58c;
mem[668] = 144'h09941daf1c14f011090cf5bae3741b49eb3b;
mem[669] = 144'hf5cdfea9103e0a2f04d9eff7f8db1e5cef01;
mem[670] = 144'h1f65f933eed6e61df59f0864e6d81f751b9c;
mem[671] = 144'h1ee0fa5a168a1f4e0ea3fd3e0a93023fef49;
mem[672] = 144'h00120c360a34ef0a17b8f8120580eceff9ac;
mem[673] = 144'h18c41159f14df1ae1cee0f29e09ce887f832;
mem[674] = 144'h1a90eebbfa44e589f8aae90aef76086510e4;
mem[675] = 144'h0145ebbb1d91109203e4e6fb19b2043ee1e0;
mem[676] = 144'hf8211f971551ef351e7109c31c2210fd124b;
mem[677] = 144'he2b3f67b1712f33a11790e9fefd118f1eaab;
mem[678] = 144'hf9f8f9481f4f11dc1429087cf232ebbbe759;
mem[679] = 144'h0fe9eca8fe800559f5baecf518ade4c810df;
mem[680] = 144'hf490fa52e9c901290297fc32e453ec7104d3;
mem[681] = 144'hf741ee56079817721fb7063ee6591f68e06e;
mem[682] = 144'he8130d9fe9f0ef5318381c831ca3f6cd1f21;
mem[683] = 144'h0d32eb0f1f430ecce1ed1243181f181b1440;
mem[684] = 144'h17fb1606ed5f031ff99012d118590153e308;
mem[685] = 144'h013be5b4ec97fbf0e91fec77f93b1c121085;
mem[686] = 144'hebd30e93f64204caeed0f9431d6c1cbeeaba;
mem[687] = 144'hfad4fb01f582e82e11090253e634e8ee0014;
mem[688] = 144'h171ae935ed81eed8054de8ddef1ce4e2e547;
mem[689] = 144'h1b0a1a9c050b0710ecbd0508f12f0de0fd18;
mem[690] = 144'hfbb9f6f216990779f7261cdc1a6a175515e2;
mem[691] = 144'h06f3ee6c0b441371e0110892ee1609d902d2;
mem[692] = 144'hf9eb0e9d0e98f746ea531f9910d0f02fe338;
mem[693] = 144'he5c518b5f9efe3391163ebb9161a13bbfcd2;
mem[694] = 144'h03641bf619a518d408410bc7e6c11a7fe8f7;
mem[695] = 144'h16f9158efa8a00ee132b1560f110e53a185d;
mem[696] = 144'hf82dff641cc8e6f8fc1312eae5abfe4d16a2;
mem[697] = 144'h0690ee7df18914551d4ce353f921e14de43e;
mem[698] = 144'he6f4e3f11aa2f854f93e1f04fe631085f011;
mem[699] = 144'h1af9fc661c30f83f037de986f559088006fa;
mem[700] = 144'hff2fe5ebe6371cdce0edf8570750efd8f4b1;
mem[701] = 144'hf4f51661f3cd0128edf8e86cebb9ffd4fb8e;
mem[702] = 144'h138ffe0cee78f41c0e94faae15be0d861afe;
mem[703] = 144'he46eeb3c0e89ed730dbbfc3ae2ddf087fc15;
mem[704] = 144'h1afa0523ef130dd8fb02e18e1f1c0e3c0ddb;
mem[705] = 144'he1a5fa381a3b1bf7f729f6b7f57de1660886;
mem[706] = 144'hf28be899fb76eb1ff268187d14d8e1580fce;
mem[707] = 144'h0e82fa580d301379e81ee52bf82909b601d9;
mem[708] = 144'h0bfe005f11a80c0a12da0dae1dd00af21433;
mem[709] = 144'hf443feeb1ce2f58216b2e6d2e4961498f224;
mem[710] = 144'h0c53e5b512d00b72e84212ee01a6e86f0df9;
mem[711] = 144'he3f0f32014f9f66def39f4b1e6b207e80318;
mem[712] = 144'heef7043702f3e6f1f96e1b9a0e1fe654161c;
mem[713] = 144'h0afe11c6e0c806f007f5072e1969f946e510;
mem[714] = 144'hfb7ae2e5f7eeedc00b9cfa24fccce877e23f;
mem[715] = 144'hf9e4e281f74ef4cf021505930fabfa63ecef;
mem[716] = 144'hebe818bc0405fa0ef6b3f189e02efad3f576;
mem[717] = 144'hea8305eae9720add06ba08e0f6a404cc066b;
mem[718] = 144'hedc009a7145c18a4f7c514a40ae1fdffeadd;
mem[719] = 144'h1187e767f683fa89e254190615ac158d1ed8;
mem[720] = 144'he90a003b08d00b5de7d1114d1513e574093c;
mem[721] = 144'he499e2ec13491117f75fe4e7e5e9e69606e8;
mem[722] = 144'h08711fe91b3e09b11445fbfffc74e4eb1c73;
mem[723] = 144'he009e10b1d500622edbdfa5dfb250cf317eb;
mem[724] = 144'hf9ece32210dde2801b2ae68dff89e871177c;
mem[725] = 144'h1fdced8ffdfa173102b1fd291426173d0322;
mem[726] = 144'h15a7f8c6e536edbe0244f81803dbe306f50e;
mem[727] = 144'h070909360191ead1ec0d18cef4ccfa6bfccf;
mem[728] = 144'h1c0714ce15d9ed02ee84fc3bfa741ce21280;
mem[729] = 144'hedf31f8c1d21045df6aef004e9da03ea1943;
mem[730] = 144'hfd4f1b8bff5e04b209f71cd211ee03c017a0;
mem[731] = 144'he5c6e95d101ee12c127ff115e713fd9f1b9f;
mem[732] = 144'hf65f009aeab8e5c0f82218051dc6f9c6fdba;
mem[733] = 144'hfd230e1909a3f746e87aeb90f34f00a002b5;
mem[734] = 144'h100e0716f898fed61c0c1b8cf5cc13591c35;
mem[735] = 144'hf90c15dae76514ce0f2c1ddcff46e99509d6;
mem[736] = 144'h17e6e717061ee7d1e80efa08e82d0a091046;
mem[737] = 144'hfed70972f616f370ec15f4821cf7142fe607;
mem[738] = 144'hf2e800ddf7e1ffebfcd515701edaf81c1add;
mem[739] = 144'headd100b1c27f4cd14ea0d9b1e40f345ec02;
mem[740] = 144'h037ce6ede3a80c14fdd8fca003841c51ec9a;
mem[741] = 144'h0795f4540d44e9b8060aec66189af59e1e2c;
mem[742] = 144'hfdba0e851b66ec971cbbe2ee145c0aa60b63;
mem[743] = 144'hfa8dfec3fe7b096c17e2e873019dfacb1bdb;
mem[744] = 144'hea9000d915270d1df4c6ea300144f785e99c;
mem[745] = 144'he9a502fa0c7b00721bfaf6bf10de040ff329;
mem[746] = 144'h15cee067198c1e86f1f40627ff35f7cd06b8;
mem[747] = 144'hee690c7ce1620657ec2fe5d01cb7e133ea50;
mem[748] = 144'hfbd11ae40f49f1c60e8d1f300941ede10369;
mem[749] = 144'hefc2eff6edfc0ce60f45e93be6351cb70e05;
mem[750] = 144'he0520de91223f5a613f40d8be412e1e9ef5c;
mem[751] = 144'he3650d6aff771bb6e893f1ae1ccaec93fde8;
mem[752] = 144'h10cdfe5c19e6f4ae1a37fb21f6c0f981ec88;
mem[753] = 144'he53ee62e0ed6028bef9d0416194605defc49;
mem[754] = 144'h07cff8d20cb0f23513a0f4cf0502e98cee47;
mem[755] = 144'hfda7e3fa155c0fe5f8cfe66deb54e5781b9d;
mem[756] = 144'h079216ee0708f0b107450c5709befc7406e0;
mem[757] = 144'h105f198eff67f3d0f0d7f7cef7b2e40de986;
mem[758] = 144'heb950fc40398fa47e4fee6970c47e82de683;
mem[759] = 144'hfa80e3ec1717e9a7e0b01d0ceb950292e557;
mem[760] = 144'h082bed1bf90b0c080934132af14b16d6076f;
mem[761] = 144'he7e2e691e9b0175ce8dce1781e96fe0be77c;
mem[762] = 144'h19c0f8e5f016e8d414f9f5f3e7c0fcbdfebe;
mem[763] = 144'h1678060717bff56a0031016fee49e3cbf53b;
mem[764] = 144'h06b3ec9d1d1ef577e2be1dbcff4a08bc174f;
mem[765] = 144'h12bf0335ef59ee3000a1feb303cde273027b;
mem[766] = 144'hefff163bf7dbf935e09f07deff31038bffb0;
mem[767] = 144'h0273e6560e23f27e12390fdce6fa04cd1735;
mem[768] = 144'hed2009511aacfe0ee702f656e0a5f1f4f0ed;
mem[769] = 144'h14f3fb9ff7680319006205d61cc1f06512c8;
mem[770] = 144'he30beffe05ac15281292f787ef01e22f00a0;
mem[771] = 144'hf729fba1e9effe7ff45b13d61877088a1e7d;
mem[772] = 144'hfab81a9f198116d2fa45f54f1e48f6e91fca;
mem[773] = 144'hf1ace072f76701faffbaebc31339f1141793;
mem[774] = 144'h1e51eb19f2b31116fbf302980d51ee0903d5;
mem[775] = 144'hf7e0feeee85de87a1403eeca02a0e4caf78e;
mem[776] = 144'he8f8ff3cf0d616410e6beeb90e531eaaeb43;
mem[777] = 144'hf07ae398089b0b05f17c0566ea02fc63e98d;
mem[778] = 144'h08fcfdf60609e6f517ef1e481393fdddf932;
mem[779] = 144'h069cfff50f1aefb8108b0c26f031e6a8e006;
mem[780] = 144'h04f10e08ee5f04161a8c0e26eb70f1adee94;
mem[781] = 144'h1d52f68aea541a9ef7dce3d8eb63eb6f10a8;
mem[782] = 144'hfb56e7fafaca09d716c30605ee7817541667;
mem[783] = 144'h012eff3bec0df203ff38ed7a0586122ffec1;
mem[784] = 144'he017f3defd4fecc2ec95192d06c301f9e41c;
mem[785] = 144'h1d41f8e802b209da0ec6e5f3eb6fe10a1302;
mem[786] = 144'h1fa8f758e6751460f21c12df13e11210126a;
mem[787] = 144'h1cef02bd152600fff0c108d20348f10df533;
mem[788] = 144'h16120afc010802f41e081afe19d7eadee2b6;
mem[789] = 144'h022deb21074802841f7318c113e2e5edff42;
mem[790] = 144'hf032f733e0ce12591207165cebc10a37e7dc;
mem[791] = 144'hef8708d7e7f9e6a6fdc0e374f2c20481e21f;
mem[792] = 144'hea04e24911830786e1ade1eb179bf3a9fda9;
mem[793] = 144'he23aee7eed14f278f133e59c19f1ece7109f;
mem[794] = 144'h11d0f238144f065ef280fcecec12eb821d75;
mem[795] = 144'he32b0f340bfd16e3e37403f40e390ba61ce9;
mem[796] = 144'h00680b2cf252077c1b770417f8e40ca7028c;
mem[797] = 144'hfe771cdd1ea3103ee3641080e8a409d71d7d;
mem[798] = 144'h14021e550d5cf0bb034f08cf1c46fa05f433;
mem[799] = 144'hed091fd5f24cfa44eacc0066f091069a1fb1;
mem[800] = 144'h1c92f42afde50e0bff8a02e91673196b029d;
mem[801] = 144'h1cc31ba603edf2b4fbc6070aef621790f088;
mem[802] = 144'hed3cf98afa651c0be45fe65bfce2f4f20170;
mem[803] = 144'h1ba9070dfdb4febaf2fa197af493193b07eb;
mem[804] = 144'h034cfd970065fd7909ce087be19afff1e8e2;
mem[805] = 144'he167112209d212d9e89deda9eb6c0af405d1;
mem[806] = 144'hfd780a49fac50660ea72019df42ff481f00f;
mem[807] = 144'h007df8a6e8751485f95c06001dc2152ee2f2;
mem[808] = 144'h1722e1f715531273f6900f40eb46159de2d4;
mem[809] = 144'h165df3cf1be819f90adc0ae3f6b1ec8efa0e;
mem[810] = 144'hec7d1699e742fdd9f9c1f25ffc23f68fe212;
mem[811] = 144'h0f37f34a060e0ecef226016c123a112aff8e;
mem[812] = 144'hefed0b8aefa2192b039a02800711f3970181;
mem[813] = 144'heb07e6980d9be1771d97fe2becf2ec21045b;
mem[814] = 144'h1571ed5e1f5b1d9ce516eb960a350e79e370;
mem[815] = 144'he39eecb0176e147b1d52ff08f922e9d90ddc;
mem[816] = 144'h104ee947eaf4e15c1eb9fbd5f7990ef40204;
mem[817] = 144'h0c750e9e1d8bf835f96115c2085fef4a13f3;
mem[818] = 144'h06df1b491b2ee005e3841ceaefff14520783;
mem[819] = 144'h1d51fbebf31efb23fb6707cc1997f33801bb;
mem[820] = 144'h140b1d87f05ce9c5115f1ba904c2fcf0ee45;
mem[821] = 144'h14b4eb3dedb2e3e4f52a02bd0c6f1c79e038;
mem[822] = 144'he243082d1ff7ea3e0c571a27ea5b0029047e;
mem[823] = 144'h1e99f0c409c6e6d8fa9719f6f678f2f608ff;
mem[824] = 144'heca405c5f13c0826f7c5f4f2f955e2f41601;
mem[825] = 144'h0e9013fbee8ee3cee4a8047f0c3f168b082e;
mem[826] = 144'h0bc1fd3202491a111413f92d007a1546f82e;
mem[827] = 144'h04f8f60e0a7ef857fc9cf3b0e3e6ec741e99;
mem[828] = 144'h0229e261feeceb16fb62017e09bb11ceeb94;
mem[829] = 144'h0c84e7acf8ecf836e2d40c30e0bbe5a8f934;
mem[830] = 144'he8cde3150baa129a0e131ea1f8abe0c60764;
mem[831] = 144'hf122055114dcfefd046b02871ce6f1e6f525;
mem[832] = 144'h19aa13c4eb3cef3bf19ff97a1d151881f28a;
mem[833] = 144'h0f610afde86912c7f370fbb804951e111d34;
mem[834] = 144'hf640ffb6e38e08fc08cde0181d26eb1d03ba;
mem[835] = 144'hed38e530017eeb44ec50fa8902b20dc4fd62;
mem[836] = 144'hf42fe51d1e2ff05ffa92fb420eaee43d0550;
mem[837] = 144'hef6c007a03c215efe0f8ea940a4e0a06ff13;
mem[838] = 144'he88d0e710b1bec02fbd2e5bf0f910257e092;
mem[839] = 144'hfd4e06e61e9bf710f388150efbbe093800a7;
mem[840] = 144'h1d7eed480fd5e768e792e5e4f9c217960240;
mem[841] = 144'hfa6d16c7e9ac01d3eab21adee4a50c3ce4df;
mem[842] = 144'h0d88ecf014860c10e3321ef4000de0d70cd7;
mem[843] = 144'hf9010bfb02e6fd9a0c58fe811de8e35202e7;
mem[844] = 144'h117713cdecf213661ab1f9a8169c146aebee;
mem[845] = 144'hf406006ee5170f981c24f2b316b6fc90e68b;
mem[846] = 144'hf3c1188216e8e6660746fd1dee92f10e04bf;
mem[847] = 144'h1ad6f9ff194dfe2c1f5de9ea0e8ef0900a9b;
mem[848] = 144'he124f7e6152ce35a10eef936f8260a530119;
mem[849] = 144'hf35de8c60b90ff73fc1e0228139a017018c2;
mem[850] = 144'h0def06fdf894e079fb27f2e8e9210b460ec9;
mem[851] = 144'hea39f22c1539f1f504520972fda0f524f6f3;
mem[852] = 144'h1700f8b30531f911e98af33be9b518d30af3;
mem[853] = 144'h09bcf2ce1d341b9613ddfcb01f5dfaa60ed0;
mem[854] = 144'he52c0afc032d16fc146e17380439fd3ffdf7;
mem[855] = 144'h1e7cfaaf05ac1080fe9f1b2d1615e8d203f4;
mem[856] = 144'hf74c06e4076feec0eb0deedc0172f57b1b07;
mem[857] = 144'he959e93c1f2200870176f167f6def83f0d53;
mem[858] = 144'h107815620911e109e62fe7c8080309a3ed6f;
mem[859] = 144'h1725e23104c2e829e70e16140188042409c5;
mem[860] = 144'h0344f545f4e3e4cc1ed3ea34febdf9aa1f9b;
mem[861] = 144'hf59ef7b8e8b70131ea6de78406e7f3770df3;
mem[862] = 144'h1e5be55efe9e03a31beefb82fa3c0ed7eb9c;
mem[863] = 144'h15e8ef11ea20f5c5e3ab199b13b91926eb0e;
mem[864] = 144'h01a2065be91f0aa0fab2133aeb2dfa5d1524;
mem[865] = 144'h0b5017ba06f01bf9e8a4f037e838f8baebec;
mem[866] = 144'he1cbe04fef67e6d019f4e31a00ce180ae40f;
mem[867] = 144'h0498e4b00281182c0a17ff5013b6f75af565;
mem[868] = 144'hede9e10d1dfa1dbcffa318e6e32b1a190e49;
mem[869] = 144'h08c3183118ab10980e91151df8c6ef7602b3;
mem[870] = 144'h1321e38c11c300fb03c717d2106c01a2f350;
mem[871] = 144'he307f797fabc178ff3abfa7bf6211660f207;
mem[872] = 144'he0a6e6c9fa08f419fc53e3e4eb79f37f0ed8;
mem[873] = 144'h0397edf41db8ff3bed4814501720ec2e19bd;
mem[874] = 144'h12c0e02504ecebc9f434f9721b451ee10227;
mem[875] = 144'h1f1afc8c19ef07121ce0196e18ae05b9f226;
mem[876] = 144'h0f58e2e2e9a5e242e70f1703031907a9178a;
mem[877] = 144'hebe1e6b70e6c035a203f0e3ae255fef4e9a2;
mem[878] = 144'h0cf0e763e36dfaad0d4b0d831a0ff085eb84;
mem[879] = 144'h0145fa2a0a31080b153cf03ffb73e01a0044;
mem[880] = 144'h153de90b14860d450e00e33efc80f43116c1;
mem[881] = 144'h19bde3b300ce0fe6ebcb1c64056c1359e76e;
mem[882] = 144'he447059dee94e6d6fab5fc561e341075ff8a;
mem[883] = 144'h05f20eb7f0a117ed0be1e600f71805e9e552;
mem[884] = 144'he76205e2e2a7013e1651e11d023c12170049;
mem[885] = 144'hea2e14b21e26e7931344fe3a0ebcf6691f0f;
mem[886] = 144'heb22f2c2f465fe0412431826f20a0406f055;
mem[887] = 144'h0350e335e093e4e9f35903fe09b214bf0b70;
mem[888] = 144'h169aef3f09edf409edba1323fa8b193bf92a;
mem[889] = 144'h13a6e1b3170f16620a96e891fcc5f051f032;
mem[890] = 144'h0b0a16970b64131319d00df9e08cf134f70a;
mem[891] = 144'h1f3ff8f7e2c20783e794ed4bff461b8216f4;
mem[892] = 144'h1ca7e507fd8d0a360cf2e00fe0d0ee39093b;
mem[893] = 144'h1d11ee79e3bef1dae6670f99e501f62df0a8;
mem[894] = 144'h1278edf90423f104e3d3e1c7fe3dee9b17f1;
mem[895] = 144'h10741e27fec3e3b111e31c1c0043f7e5e686;
mem[896] = 144'h09e912830b58e4d31613e8a4e9f0f9261b81;
mem[897] = 144'he1f7f129f60e051c03881711ec3a1946f0fe;
mem[898] = 144'h1b5511c2f6dbf77fe9dc128d097eeeb2eeb7;
mem[899] = 144'h0cb6f627f6a6ff55f6a308c91e2519ecf8fa;
mem[900] = 144'he57f045eec12e7bd0b61e97ae28dfe340942;
mem[901] = 144'h10721fea086ce810f99c184ae4e00cc10017;
mem[902] = 144'hf4b3fef90c11e056f123e4bde5f4f8530138;
mem[903] = 144'h1802004e1955044315220a5901c1102b081e;
mem[904] = 144'h16241589fd3c1aeaf715fca8e0470136074a;
mem[905] = 144'hf73ff58cfba718901d03e6d6e6b7f2f8199e;
mem[906] = 144'he7a8fe051dd8190304de0e0c1ee90acd0da4;
mem[907] = 144'h13630d8ef3bb023df911091d1aede5eee735;
mem[908] = 144'h12ec075709f9f379ea2f04711f36f03403f3;
mem[909] = 144'hee8404ee063608f114c2f48b14a9f7bb0cc8;
mem[910] = 144'h04e415cdeee6fd7fe07bf653ee55eecf099d;
mem[911] = 144'h1fdf13bb079e14f90e4feb661491e77301d4;
mem[912] = 144'h1b790995f262e53016d5f3cceadf14e416fc;
mem[913] = 144'h02ea0c08e03cecbff0e4f666f64be3d51cf7;
mem[914] = 144'he59e0a0f1b24ef56028f1a770756f6f9f597;
mem[915] = 144'hf38e09abebe306cd1d3c1ccc0378f0e4ef42;
mem[916] = 144'he9e5e0c901441a8dfc891d63000012f4e254;
mem[917] = 144'hf4d4f788f9baf333146f09e5e443ff0fe2ea;
mem[918] = 144'hf1bcf4bcf6aa107a01cef53103ee164dff6e;
mem[919] = 144'hf2ef07701e63f621ffd1ea01e4311a4e0d3e;
mem[920] = 144'h021019f70fd3e3b50bcde3f11a5bf04506d0;
mem[921] = 144'hfdd40ad9fe6c1b9dfa711301008f193dea0b;
mem[922] = 144'h0d9a0ebae37df247eaed0bb2eca5e65de071;
mem[923] = 144'hff2ffc550ea01c74f606ef12f462eef70c6a;
mem[924] = 144'hf0adf98fe4ec0984ea4a1338e26006c9e689;
mem[925] = 144'h0ee4ff7c1dd10bdb0b9615fc0c1c182b0528;
mem[926] = 144'h11a6f0501184ecd5ea20f2cfef9fe23100d0;
mem[927] = 144'h074f09ad00affddcf78de0781664e270e746;
mem[928] = 144'hf83c102a10daf38ef1db043c062af944f976;
mem[929] = 144'h1bd41b6a0182053dfef2fe030b05e025e5f1;
mem[930] = 144'hf54601d00029f6271bf90221fe0ff73e034e;
mem[931] = 144'hf931fed2f6700defef99fe7b11421cc4ff1e;
mem[932] = 144'h135705bf0904fd39ffd00dbaed76180bec68;
mem[933] = 144'hef240070fc5af81b0c4b035802251439e712;
mem[934] = 144'he604e491e4a700df09adef59e493f673e444;
mem[935] = 144'he3fc1caf1f75eaf907981725f360fcd7075e;
mem[936] = 144'hfe4be758e69f0cc711781e57fba71c321956;
mem[937] = 144'hfcb61d10141ae9a2e2faf3ebfadf1f5d1982;
mem[938] = 144'hf7f8040b1ae7131fe5220125f6bd118c08ef;
mem[939] = 144'hf25af88dfb90ffc7f29c07d7ead51a3dfa5b;
mem[940] = 144'h1feb1d85f66ffc3d08d5e28aec6d028a07dc;
mem[941] = 144'h1786f25a16ca076d1dbdfbb6e596f8f5177c;
mem[942] = 144'h07ffe00ae9350cad0a2cee0c0a5a01b60c4f;
mem[943] = 144'hfec9ee08e0f6f60e0f49ea241505efc1f11e;
mem[944] = 144'hf2d514690a4f15ecfa94f7631f1efd2eea07;
mem[945] = 144'hfb05f8d301440285e5b8e6ae0b480f270a3b;
mem[946] = 144'h01ad14d91368effa0a4d137604faf11e0f98;
mem[947] = 144'hf58cf872ec1ce8f60fe3068e0b870f3e0cc2;
mem[948] = 144'h1dbaf70ef5cf19e6e9fef39dfe770b060ff9;
mem[949] = 144'h0d680fe2e05209ff1a9300c8f890f4f8fe0c;
mem[950] = 144'h1bd3f4ee1a56fc3ceb28150411241627fe6f;
mem[951] = 144'h06050fc61b0714fa0b20fa06ff540d11fcc5;
mem[952] = 144'he54aeb23ea3b0005f594f3430ec613641dfe;
mem[953] = 144'h0d5be31afacfe200fd95e4e711fbe5410c0d;
mem[954] = 144'heec3e1ebf31718130300e4fd1f13e076e814;
mem[955] = 144'hfe5907bf0f820f580729198118331f14f349;
mem[956] = 144'hf4811eefed9d04abee0af7effc2e0469ef51;
mem[957] = 144'he60f01cdfff9fbd3fe8817c4e98febcdf614;
mem[958] = 144'h1a71126b0336e1731aa91a52159bf642099e;
mem[959] = 144'hf05df8dc1c7fef0be528e26318bfedf11953;
mem[960] = 144'h13d1121de3fe035303eaeeb9f98008ae1c59;
mem[961] = 144'h1e380204f805ecaf1bd40e731ed7fdfce45b;
mem[962] = 144'hefc91d98f66bf8c6f94204031a53f596fa63;
mem[963] = 144'he841f4eb157c0551f8f905daed21e048e8c8;
mem[964] = 144'hec98e1a1097ef2ae0caa150009dce481f3b9;
mem[965] = 144'hf4f1f997f56d1630090ffb38f803e604ea91;
mem[966] = 144'hed2ce7cee6921e5deca6e8840d80fadb146a;
mem[967] = 144'hec3418a8eba805eaeca813530ac70b490e8f;
mem[968] = 144'hf8471b5b039600f8e126ed52e669e67504c5;
mem[969] = 144'h13b80d8be065ec8a13c11e701a94f6351dfe;
mem[970] = 144'h119f17dd05afec1c15580497feed07351192;
mem[971] = 144'hfd2be1e7e8960fac10c6ffe4fca709f9eb72;
mem[972] = 144'h13bdf52d1813f5ae02370a60ef95ee4802d7;
mem[973] = 144'he2c715aeebc014691264120c13c9e89a11df;
mem[974] = 144'h0affe343f9c6eb25f7f3026b1244093b0df1;
mem[975] = 144'he7260324f9bd0b6608eaebc1e56ef0e1102c;
mem[976] = 144'h1a7504251ca904ac0db90d3e0d6b0adc1de0;
mem[977] = 144'h1ecefa43fe1e11f5ed3ce6a7f851ee0b19cc;
mem[978] = 144'h02bff414fd5bfaf2f093100ef814e591007d;
mem[979] = 144'he590e698f896ec7b1611ee6b156a167314e5;
mem[980] = 144'h11cc1ea1f6bf120fed1a13b4e322e7f70ff0;
mem[981] = 144'h00f81ba0113f11d30a5313fd1e44153afd27;
mem[982] = 144'hfbace9350febf66cea011888e160eebe0a5c;
mem[983] = 144'hf2eefcd303f9142afa76ebba1fc5fa0d1f07;
mem[984] = 144'h018818f7fa92fcdbea3f076ee5641f22f5c1;
mem[985] = 144'hee2deed3e56a08c41dbaeefc0b5be5a9fa20;
mem[986] = 144'hfc56fc0fec85f9a0e91ff858eac0f1ab0264;
mem[987] = 144'h1b4ef6e71fcb1feff096fb54167ffb5a1045;
mem[988] = 144'h0f14e5a40373f0f3f669f8f80a69ec771821;
mem[989] = 144'h1ae6f661fd4e050d105f069e11cdfd79eb66;
mem[990] = 144'h17da070a002508ba191118f70272f4bc1232;
mem[991] = 144'hf3ca0677f89b1c70ea1af4b909431e89eaa9;
mem[992] = 144'h12ba16fe1e00f6f8f139ef55f241ed59f13c;
mem[993] = 144'he353047b19330ae8f4a113f1f3e40bdc1d67;
mem[994] = 144'h11f913031cdf08f71644e097eea4fce6e841;
mem[995] = 144'h0316f7a4e097e40ef7ce0ac7175a0c761b82;
mem[996] = 144'he1b2e876166de3940b5a1a3116effb391688;
mem[997] = 144'hfba2fb3409490cb9e0da09290d87faea076f;
mem[998] = 144'he261f7af1222eca61f20ec56ec440da2ec7d;
mem[999] = 144'hef0504f1fffff5d605fe1f00089b1a34022d;
mem[1000] = 144'h1dfb1ee0f5321561f272128b11dae747183c;
mem[1001] = 144'hf30fea16fce71003e821ebb505ab08131b0a;
mem[1002] = 144'h0dfd0dc5072d0cba19c812681d55fa1f05f6;
mem[1003] = 144'he132fc8e0329ff1df9b21bcfe989161efa26;
mem[1004] = 144'h0e4410d618941943005504e40145011e159c;
mem[1005] = 144'h1a9109dee2daf6f10e5ff8a4ec1cf86a01d3;
mem[1006] = 144'h1a7ee617180709ba1defeb29190d15da0a75;
mem[1007] = 144'he73afbda0663e671f49b015c0d11f9daea8d;
mem[1008] = 144'h09f9032def4a063ee79a125602e4eff41d07;
mem[1009] = 144'hff7b00d1f3dbe43bf84308821a431fc51d2d;
mem[1010] = 144'h0167f240e88312671c7cfe84fb1bfd19edc0;
mem[1011] = 144'hf456f828f3c7e4170d49ea05e2a803ff150a;
mem[1012] = 144'he74a033d02bdeda2e7f80924e2871217e65c;
mem[1013] = 144'h131be2b4fcacfea31745ebc4f623f072e75c;
mem[1014] = 144'h0b1a1065f680fea1f00216060b49e5f11d36;
mem[1015] = 144'h085f07d6175219b9f8ba17091158172111ea;
mem[1016] = 144'hfc040c56edbefe46fad50b001b1501811d3c;
mem[1017] = 144'h1eb40f9a1d9df3c4fa1c15ce001df01ef4f8;
mem[1018] = 144'h1e34e43e08ba09a7f9110f071e821ef9e7a3;
mem[1019] = 144'he13a11fe0ee5f9a31a69e08fe3c7f7ed0fc6;
mem[1020] = 144'he4c3f9bbf6c206f3ff1ff3170e1ef01dfd7f;
mem[1021] = 144'h19400ffe0361eb55f0db096e0ecc1516f6d7;
mem[1022] = 144'hebf3efbe171a0f2feee3f9f4f26cf99ae5af;
mem[1023] = 144'hfe39153706010cc9fa66ea8a19a106f9f6fc;
mem[1024] = 144'h00f517f2f0f30a4e1baa08eef43e0b881d22;
mem[1025] = 144'h08da052b0f48e44405cde98af1f91b341772;
mem[1026] = 144'h1ba5e0f4e480f148f821f006f183e1dcf2be;
mem[1027] = 144'h1f8efedf15921c27f61f1191075cf5a7ff0f;
mem[1028] = 144'hebf217430b1411b3061d083d08ff05b50642;
mem[1029] = 144'h02cbea2f1c34f91aec0b1fd8efa506cbe552;
mem[1030] = 144'he75d177fe14118e5f7cced0afd8be9ca1d0c;
mem[1031] = 144'he271ef56f798e772070c14bcf08bef091f76;
mem[1032] = 144'h14000ee2116c0ea9f3b8edd3eeb1e6a30f9a;
mem[1033] = 144'h0d201e32f2d2fb3e0723efc21736fb46e37c;
mem[1034] = 144'h16941c4ff13ae896e70fe2c4f38117500728;
mem[1035] = 144'hec75f4b20074e739e39b0b02f60bf0dd1875;
mem[1036] = 144'h0ab5e0261f1efaa71bdf0f28e6bf0679e9ea;
mem[1037] = 144'he676f64b1afd15f80bfd1eea15abf365f07c;
mem[1038] = 144'h19c9f99001690af90a0511e9077fedb2f830;
mem[1039] = 144'h0cfc0255e153f8edee531d6412f7f88619da;
mem[1040] = 144'h0fbb0fe307f0e54a02ff0c76f9970a5f1031;
mem[1041] = 144'h17131f1efc13040f15caec3cef160a1be7a2;
mem[1042] = 144'he96ae6060d301604e44ef3b5fc7408c6fccc;
mem[1043] = 144'h0e4d12e3f1fd014b1823eda0f178f5450a36;
mem[1044] = 144'h1b3a0baff06c0c981177e7950069fe370e1e;
mem[1045] = 144'h1ad8f7001e960326f0f0ff8e106404fae12a;
mem[1046] = 144'hfbc41682e11f03d2fecf0bc8ff6a1a101a2d;
mem[1047] = 144'hfc9ce84f19d205dbe10df9f8ecd4041d08bd;
mem[1048] = 144'h19421bae0e8af9c5fd680b7dfd1ce58c1ae0;
mem[1049] = 144'hf9bff7a6f54a0827eafbe611f77900a6087c;
mem[1050] = 144'hf3891223fd100dc2f36404990aa21bd5ff51;
mem[1051] = 144'hff611de004c6e3711b2d08b6f630e7c0066e;
mem[1052] = 144'hfb78157514931d7de47d1b1aecd5e470fad8;
mem[1053] = 144'h189c1f4a03da1e7e1c02fb9e1ca815fd0d39;
mem[1054] = 144'h0b1e13c80f55e2bc06fce343f99507a60b32;
mem[1055] = 144'h1b9ef2ae04c7e504e2d30125fa33e4d4e5f3;
mem[1056] = 144'he34713adef13128b07e50736013c064c1206;
mem[1057] = 144'he2ec1d9ff8c30617fe9eea981652108d035c;
mem[1058] = 144'hfaacf50a1ba10f64eb9f1de20829e3ceef61;
mem[1059] = 144'h049c0c411203e99c1009ead30fcae4f4fd37;
mem[1060] = 144'h032ee23de7c41a1b05181ad104efe22a0466;
mem[1061] = 144'he8ece3d3ff830615eb9800a118b61d7fe598;
mem[1062] = 144'h1526e8acf5c5eff2f37fee05f6a1048df87b;
mem[1063] = 144'hed9df03a0762094d0113e464ef4a0010f17f;
mem[1064] = 144'h150a0dfa15e0e76df562e6a9ed4303ba0b22;
mem[1065] = 144'hf8270a060e2107ec0b8f1f5605b0f1ccec92;
mem[1066] = 144'h1c691cd7111d19af1b88f4bbe9ecf35df83c;
mem[1067] = 144'he3f2f86de40ef6e0e35ef304e3c61fb2009d;
mem[1068] = 144'h0fc5f2ed1719f27018661e9b1c9c08740b78;
mem[1069] = 144'hec8306af00050c16e5e51825ee541c921102;
mem[1070] = 144'h0bfc0dab07de1f9e11781e8602fcf952eedd;
mem[1071] = 144'h1beaee72e5c214eb1b4d1144eb5d05211f28;
mem[1072] = 144'he4c5fe551132eac4e29de9d20665f77704a8;
mem[1073] = 144'he3cdf2d10e2d0e0802be1661ff9701e2103d;
mem[1074] = 144'hf1f0f38ee6f814df04d9ed5d0238ead4f0d9;
mem[1075] = 144'h0de7166302040962fbce0e73ff39fd55fac8;
mem[1076] = 144'he1fffc2ce29906f80bc607ef1842eb86ef0c;
mem[1077] = 144'h19b215fafc45e3d1028b10e8f62ee40efa81;
mem[1078] = 144'he632173f0e1cf0f50d88e42507280bab0913;
mem[1079] = 144'hf8d2eede116ae3df02970716013a1ca50699;
mem[1080] = 144'hff5dfe7de9bff8fae92d0c6ee6d71ac61c00;
mem[1081] = 144'hf53f0b9fe93305a4ffe0fd3de3c80273e1a9;
mem[1082] = 144'h1c3cf7e514040964e67afacbfb74f988e0bb;
mem[1083] = 144'hee44e0d21ad9085510b1f1d6ef9cf4a108f0;
mem[1084] = 144'hf40efadeeada191f0384e1a41cc2e8b5f60e;
mem[1085] = 144'h09b6e0440d58011804a0e68106fde041061c;
mem[1086] = 144'h09e21083063cf322fbde19d8fe1eeeeae905;
mem[1087] = 144'hffc60042f4700cfcfbf8e6b305db08d916e9;
mem[1088] = 144'hf0fc1fbae90e00681076f0fae79e0316e0ff;
mem[1089] = 144'h1014e1480671fdb31d92f6e81778f5cae8d8;
mem[1090] = 144'hf0f4e5d2faafeb89f904e60bf9490765fe7a;
mem[1091] = 144'hec0d136807d41ef8ff8210f41bcbef26e4fc;
mem[1092] = 144'h10ecf6c5fe1de6da101ff7d8ec600b711e46;
mem[1093] = 144'h0d91102a04001867ecf601531b2eef3ef862;
mem[1094] = 144'hf74710eafc1ae05afffe1d0dfa80f4fcf186;
mem[1095] = 144'h1051f058e7f90a0e0c55079d0b2f1c600eda;
mem[1096] = 144'he6071386eb20ff54f0db015c171f02431944;
mem[1097] = 144'hfc9bf9ff0a23e61c177bff3ceb04199cf2f7;
mem[1098] = 144'hf2ccea6f12e0f7451b910391eac10f1714c4;
mem[1099] = 144'hfad0ea3a029312ac14a31a3efcaa01471bf0;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule