`timescale 1ns/1ns

module wt_mem1 #(parameter ADDR_WIDTH = 11, DATA_WIDTH = 144, DEPTH = 1100) (
input wire clk,
input wire [ADDR_WIDTH-1:0] addr_a, 
input wire [ADDR_WIDTH-1:0] addr_b, 
output reg [DATA_WIDTH-1:0] q_a,
output reg [DATA_WIDTH-1:0] q_b
);

reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

initial begin
mem[0] = 144'h0ca90cd4f396f2d8fd8efc400cf807a30bee;
mem[1] = 144'h0a5e0cf807d60211f83ffb66006b06c900f9;
mem[2] = 144'h0e15fab2f383ff940cad08deff7bfb92fc49;
mem[3] = 144'h0f32f822f84dfdf3fcf50339f37102e606aa;
mem[4] = 144'h0687f1aaf220ffbf059b0078fed0f12ff2e3;
mem[5] = 144'h0b1ff5dff3ae0450fd7b02b3fbc7ff39f6fe;
mem[6] = 144'hf6a2fab0f02504ec08b103290aa60545fc2a;
mem[7] = 144'h0679f6adf1e0004af31efce50f74f340fe38;
mem[8] = 144'hfcd3090af28707cbfa0cf35a0a3d00e9f41a;
mem[9] = 144'hffc2f3ac0b9700fcff7df85ffe0f0b20f685;
mem[10] = 144'hfee707c8f5bc0d2e078a031cf34f01faf99b;
mem[11] = 144'hf426f3a504c3071a046407def386fa8502a9;
mem[12] = 144'h04eaf36af413070d0428f2f300f8f409f469;
mem[13] = 144'hfecd0a570517f6b4f56b0c64f315f5270055;
mem[14] = 144'h0e6cf6fc044bf834fbd2f5a20d36f291f139;
mem[15] = 144'h0faafae4fcfffb1d0c42f6c90ecffe6ef3e3;
mem[16] = 144'hfa4a0186fb6301a5fa5707fa0f3e038afd2d;
mem[17] = 144'hfb2101aef1ce079505d1f97109650c44f13e;
mem[18] = 144'h07c60f4bfe9afce00b69f80e0eadfc340921;
mem[19] = 144'h0b1b0f70fa6d0eaf0167fdef01d20062fffd;
mem[20] = 144'hf4c20a910ba1f0650394f314fdaa00740d07;
mem[21] = 144'hf4680e00fc0e02f9f6fc00c90c9aff4cf874;
mem[22] = 144'h04c5fb13f63cf3dff2c705410003f484fd7f;
mem[23] = 144'h0ba3074109e40d30f748fcd5063e02350f5f;
mem[24] = 144'hfcd107ca08d8f97a0f55f629f814f5a30fcc;
mem[25] = 144'h0ab30bb309dc034208870c98fb97fe5ffdc7;
mem[26] = 144'hfcb3fb7f0e320c54f6a6f39701aafe32fec5;
mem[27] = 144'h096b055cfbf00186f73600d8f884feac0f73;
mem[28] = 144'h0db00940081fefd6f7050a0a03210d4501e1;
mem[29] = 144'h0b2c0f3f06e7fc7b0189ff2c03e50d7a0409;
mem[30] = 144'hff09fe7b07880f0cfab3000b09b0f1f0f635;
mem[31] = 144'h05db07def4090d2af855f3ce0d5c0619f5f4;
mem[32] = 144'hf441f994fe0fff430888f8ff052f0216086f;
mem[33] = 144'h00b2065ef99e0ff3fd890a09ffedf170fb74;
mem[34] = 144'hf7e1fcdb02b5fd99f5d4fbfc06450b60f721;
mem[35] = 144'h0609ff05f8e003dc0e60fe50fe37f2b102cf;
mem[36] = 144'h014309b409a20da202d5f1a8f9b208bbf90e;
mem[37] = 144'hfd51fc31fa99fbe5f0bb0f4ff63dfeab01d7;
mem[38] = 144'hfb81f7270c250b3602b90d59fd42ff2609cb;
mem[39] = 144'hf908fc0bf315f25d08650c670a29f5700b8b;
mem[40] = 144'heff305b9f7c5fbf3fbf5023a0ca8041e0f73;
mem[41] = 144'hf843fedff62b0bfbf2cf00e9098301d5fb30;
mem[42] = 144'h0bf3007bfdfa0366f1820151f66a0b7001ee;
mem[43] = 144'h0c9df9daf415ff4cf18ffb2efe1607e9fc74;
mem[44] = 144'h0ad1ef8800b2fabf09650b80f8e7ffe406e7;
mem[45] = 144'h05f1f158f60dffdffb0109adfc35f774fc6c;
mem[46] = 144'h0d0900720d6bf9f8fe13f16f0951098805b2;
mem[47] = 144'h07920c3c06730a78f29a05f4f4e70720f355;
mem[48] = 144'h0c940fa0ffc90594f0b302a60475fcfff274;
mem[49] = 144'h0e6e03660b87fc8606b00d88024dfc5f07f3;
mem[50] = 144'hf8b4f9540b990065048ef6b2f7b90c4efccb;
mem[51] = 144'hf9fc0ad204befc010590f6e1092afd2503ba;
mem[52] = 144'hf5340972f1c8fa69f6bcfd560ecd0fbdfcca;
mem[53] = 144'hfbc9089bff24ff26fbf20711fad706750dbb;
mem[54] = 144'h0eec0b7c050bf9650ca10e0500a8f5f80f09;
mem[55] = 144'h07b3f2baf105fdfb097701b7f19604ee06df;
mem[56] = 144'h0a8b05e90ec7f447f0def34c0753ff6f078b;
mem[57] = 144'h03b7f53c0cb8f1ccf7320919fbd2f16ffba9;
mem[58] = 144'h03a802dafab1fe4102ddff74f0100450060a;
mem[59] = 144'heff30015efe8f4bbfc0309ce00d5f9910418;
mem[60] = 144'hf33d0c3b07f400f60545098ff5140b0a0427;
mem[61] = 144'h0afcfe730f35f850facb0385003c0aa9f589;
mem[62] = 144'hf352f6b60df2f8daf0f1f8560890fdf60238;
mem[63] = 144'h054ff16e092c0b2ef9d7f92cffed047fffe2;
mem[64] = 144'h0a9cfaef07b3f6280589004d0a6ff1b20e82;
mem[65] = 144'hfd9ff8b6fe3a0420fce1f3160aa001c1081a;
mem[66] = 144'hf47ff437fabf0748f8f7fee70322f09204d5;
mem[67] = 144'h07b60558f49efa790472f9bd0f360051f4ca;
mem[68] = 144'hfc3cf147f490f279f517023b0c0cfe130c6a;
mem[69] = 144'hf5eb0c88f1e20a7a08a00858f8ca0c650960;
mem[70] = 144'h0a6afecb0d5df1a9005003cb08fa02d10caa;
mem[71] = 144'hf59e055d066b0cde034dff00f0f7f7f30762;
mem[72] = 144'h03ecf248025ffd01f33d0f06086802bc0a0f;
mem[73] = 144'hffedfe790f04f95bf5af065f0768f3f60816;
mem[74] = 144'hf7900f63012c0f70f80ff038feab0239f41c;
mem[75] = 144'h092f0819f16d0a5ffd51f1e3f0c9fe1d050c;
mem[76] = 144'hfd9a0f33f84103f70b140cca0b9bf4adf9cf;
mem[77] = 144'hfdd7facb072cf2b0f5f9f40df6cd0f840de3;
mem[78] = 144'h0f2b053bf145f1ee0b86089202010e7b0424;
mem[79] = 144'h028ef609f1a90e8cfb9f0d24f8dc0ef6f378;
mem[80] = 144'h00bf0fbbfffaf5c20201fdbf0b86f17e0f4f;
mem[81] = 144'hfe700be10faff169f04dfc0bf49df99cfadb;
mem[82] = 144'hf289f20c0e8104d4f84df98af12af530f4ac;
mem[83] = 144'hf358ff770dcb03adf80e04cafda90b5c00ce;
mem[84] = 144'hfe530b9800eb00d3f68303780e680883081a;
mem[85] = 144'h00d603280b140c2509df05530e32f1def3db;
mem[86] = 144'h0da00b70f61df0e8f15bf03efcdb02c8ff28;
mem[87] = 144'hfdd30a10fa560d09fb5604920e28f68e0f27;
mem[88] = 144'hf379087b0e4c063dfb880c47f05406d4f2fe;
mem[89] = 144'h028ffb5605330afbfa84fe10015b0eec0a67;
mem[90] = 144'h04bafa9d07b809dd083df83a090cf09efdd4;
mem[91] = 144'hfee8f566f874fd95fb9b0fdafed303acf6cd;
mem[92] = 144'h04e00612fb4cfe20fd72f9b5f458f51407c2;
mem[93] = 144'h0db0f0edf7ac05e0fc2900ebf2a605a8f408;
mem[94] = 144'h0b0af9ca03bdf51bf014047c0beb0820fbb3;
mem[95] = 144'hf7c90051f4d10c5b02fb07d7f960febf0d20;
mem[96] = 144'h061a03810691fc38f08e0f4802adfa8aff47;
mem[97] = 144'hf813f511f4e0f960f4eafb1a038b0baa07e4;
mem[98] = 144'h0bd4f288080405440177f432f209fe330634;
mem[99] = 144'h0091fa7ffd8002ebfd53f9150d1ffeabf910;
mem[100] = 144'hfb83fafaf01df16df4cdfb7fff730ffe09aa;
mem[101] = 144'hfc36ffad0ecff1b8fa2c00fcf210f65b0a78;
mem[102] = 144'h0a3d0ba103190d940929f71804790d53f1d4;
mem[103] = 144'hf3020e08f031f718f62602fafe84093d0951;
mem[104] = 144'hf079ff6df14df6c500950792fafef39400e2;
mem[105] = 144'hf3e3fd11f4d60f2af817f0a3019ef7b1057a;
mem[106] = 144'hf5d4fd610f97042bf7a90ccafdbfff790e7f;
mem[107] = 144'h0c800ab30cea052f054f032507caf2c70553;
mem[108] = 144'hf5a4f8c9fc29f625f154fd24077b03660b09;
mem[109] = 144'hf9170693f663f56b00360ae8fe9905a60efb;
mem[110] = 144'hfa02fa9803390d3ff570055d05790e830343;
mem[111] = 144'h0ae906dcfd12fe480f63fb440712f5d502ee;
mem[112] = 144'h062eff1ff3b30f960699f9ec0c7e0661fe30;
mem[113] = 144'h0ace038c05b3f424024bfaaa0054049e074f;
mem[114] = 144'hfd740410faaf0e0a0151f96efa5508890405;
mem[115] = 144'h0af8f82df1cd0603f574f82b0cb4f86606dc;
mem[116] = 144'hf49ff397fd9a097d0ea5fac3fddaf83dfe1f;
mem[117] = 144'h0b010a3cf99af7d3f01f0cd60172f29607df;
mem[118] = 144'hf395001c09affbda075ef229035ef1e7fd19;
mem[119] = 144'hf967035404c3fa84f6e0f41e0938febdfe87;
mem[120] = 144'hffa6f5590719f272f4ee0826f6e809f0f562;
mem[121] = 144'h094dfa1ff41404fe0069fa55f43500e9f6c2;
mem[122] = 144'hfa060b76f5bf07240f88fdaf0160f65efe8a;
mem[123] = 144'hfc75f87ffb3009d201490a650875f7250933;
mem[124] = 144'h0d79f61bff9af818f14204fe026301fa0f6c;
mem[125] = 144'hff7c074dfed502d5fd6d0aeef1faf0cbffc0;
mem[126] = 144'h0cc2fa6e0e9cfc65f96ff0b6035cf8e0fc33;
mem[127] = 144'hf3500285f3f80796f86b0c9ff1ebf9a80af9;
mem[128] = 144'h050ef5d7012cfe510a3af7b0fbab0a3df7ce;
mem[129] = 144'hf98009020cb4eff8f34dfafdf68e0954ff33;
mem[130] = 144'hff89fd290440011f0937f53bf2eb0592f166;
mem[131] = 144'h0acf0f1e0596f5530c4dfb750a840425077f;
mem[132] = 144'h0a2102fdf72dfa1307d4033303d50c58f267;
mem[133] = 144'h067c0a20f77f0b220d0d0524f062026f02c0;
mem[134] = 144'hf58fffecf75ef080f30d0077f0b906dcfacc;
mem[135] = 144'h0704fde0f5e4f081f1c6f7cef33df28c087a;
mem[136] = 144'hfd0df965044af770f3d40adc040cff8c045d;
mem[137] = 144'hf8630d160d26fd120214fd8905e80aac0fd6;
mem[138] = 144'h0137ff45f34af7c3fb5a00ef04e4fb70f293;
mem[139] = 144'h0e7cf921fa4e09d70cf4fba8fff90bc4f2b7;
mem[140] = 144'hfbd4003f0704094a0ccef3fc00f0f5b4f502;
mem[141] = 144'hfa9df2fcfeb4fa840ae4f1bcf5d90a67f629;
mem[142] = 144'h0f6ff9e5fb08f60eff7d0cad0b1c05acf5a3;
mem[143] = 144'h0088fb0ffe73f63af4fcfc26f65d0f33ffe3;
mem[144] = 144'h0298f3fa00a7070ffca40b77fb0a027f0860;
mem[145] = 144'hff010471fe5ff6ff06dd0b35f39a03310da1;
mem[146] = 144'hfeba046ffd4cfcc00bd3fa25f57106dd0988;
mem[147] = 144'hfc15f86ff8ef04dffae909c5f1880201fe51;
mem[148] = 144'hf5d00429051ef789f69b00d1f75ef197f4ef;
mem[149] = 144'h05cdf4840dbc0e7cf2fa0131f472fdfaf987;
mem[150] = 144'h0963f77a0b66fffa09130c6e02bbffe5f983;
mem[151] = 144'hfc39079700a5fd5708fdfa670822f1a10f1b;
mem[152] = 144'h0fcbf8c3f657f4e70b93f87cfa8005bbf4a9;
mem[153] = 144'h08e10e640d50f57df7aef89cf93305d20bc8;
mem[154] = 144'hfa390fb2018206390d65f7b10139fba703f1;
mem[155] = 144'hf69af2d70b61f0540a46083f0cf8fc980084;
mem[156] = 144'h0ab40d260bacf2c1f56b0f65030d068a0be0;
mem[157] = 144'hfea9f02dfeccfd9ef74eff17f4cbf9760300;
mem[158] = 144'h01dff7af051007c3f1a90bf00e1b0bdffa28;
mem[159] = 144'hfe1df52dfdcf0e9c03e3f1db013a084303bc;
mem[160] = 144'h0e7e011f0e9f0915f8e20f89fd020f450636;
mem[161] = 144'h0d3dfab30c90fe960a6e0bb4f7da06c3fcad;
mem[162] = 144'h00800b56027105740933f383fbdffeae0f82;
mem[163] = 144'hf8a9092708d90898f688010cfb740141f5a7;
mem[164] = 144'h0aa709010019f883054dff84066afa9cf7e9;
mem[165] = 144'hf9b003440ab8f4350b87f2a30b39f2b40283;
mem[166] = 144'hfbe80ed20c630e3106690252fd49fb7bf940;
mem[167] = 144'hfdcdf7ee0da109f7f55ef18d0eec048af808;
mem[168] = 144'h0fc5f927068606bff865fa21f6390c5c0d57;
mem[169] = 144'h0b810665f438fe58f4cdf4e80d3d00580999;
mem[170] = 144'hf349037bf68403700eac0113f12b01260a45;
mem[171] = 144'hf4f5023c00cef30af500037d06a4f6b3037b;
mem[172] = 144'h0b960a05007bf1950b5ef9730799f6db08ae;
mem[173] = 144'hf03f0643feb5001b01740d33f599f492088b;
mem[174] = 144'hf075f715f071fe49f40af9a9f4e4f1faf764;
mem[175] = 144'h0398059cf90fffb1f9d1f87effc7fd9ffe94;
mem[176] = 144'hf8390c60f5b9f5f8fa57f088ff140a1b003c;
mem[177] = 144'h0e220024f75ef0d705040bf8f35b0c26f018;
mem[178] = 144'hf87e08380eacfe130edf0a83f1420d6afdee;
mem[179] = 144'hf3cbffcb0ebbfca7094402acf976fc5ef438;
mem[180] = 144'hfd0007910333f48cf70504fb0f640758f289;
mem[181] = 144'hf074094408c7f9640e6af0c5046e088d0249;
mem[182] = 144'h0c59f474f8270daffc3603caf1000f660ef1;
mem[183] = 144'hf026fccefef60abcf63b06d6f2bff3cb0d16;
mem[184] = 144'hf94c0e190c5b0fc0fa500e9d0b5405f80801;
mem[185] = 144'h09d3f2e4f16a0cc60b270949f3effcd4ffdf;
mem[186] = 144'h081df9ab0287f0540e39fd8cf7ac088b048a;
mem[187] = 144'h061cf7b8f2440b64f9820b66f3e802f5076f;
mem[188] = 144'h0c2205bf0deafb38f7130144058df7b90641;
mem[189] = 144'h0a11ffea0570fd0801a1f8b709aaf8d1018d;
mem[190] = 144'h0443f6fff9800d260025fdcbf0f9fffb0fe6;
mem[191] = 144'h0b8f0bf3f997f5c909860ec101d7f4df0a45;
mem[192] = 144'hf059ffc6011afcaf08b2f4c70e4efd18fd67;
mem[193] = 144'hfcb1f8390ad00badf817f7e90ff40011ff51;
mem[194] = 144'hf7660f3b03b5f440f5c30f1706b20fa4fb08;
mem[195] = 144'h0608fa2f0602fcaef0c3f7630413fd59f8af;
mem[196] = 144'hfd7c0954f667f633fe60f139f53bfff50b4d;
mem[197] = 144'hfa3f07ce0039f1a10ba00e970a660760f686;
mem[198] = 144'h03e5f3bc09a7f1a50cd9f47504e00e62024d;
mem[199] = 144'hf571090f0bb5f294f2060933fbedffddfaa8;
mem[200] = 144'h0026fcfcf248fc83f8e4fa6e06cff0300dad;
mem[201] = 144'hfaca09bcf8280093f8a50161080df48b00ce;
mem[202] = 144'h0b6306df0be10f3e0346053c04820c67f4a1;
mem[203] = 144'hf68a0be70fe2f190f4f30d8cf2150418025f;
mem[204] = 144'h02030b3c069ff2c2fff4f0610ba3fc4cffdb;
mem[205] = 144'h0e1ff7a7f75df97c0e8f098507ccfa8ff56d;
mem[206] = 144'h0a31ffb5fa2cf64ef9b50d23ffbbf73907ed;
mem[207] = 144'h096ef813f9e10c8305b0fd57f283fada0612;
mem[208] = 144'h056efbb40ad5f153f0e0fb240def0848f223;
mem[209] = 144'h04b2fc32f1bbf2730fd9fe62fe8afe65055c;
mem[210] = 144'h0cbf08eaf4c9fe0c0dc5f6f804550dc6f188;
mem[211] = 144'h01b403a9ffc60624f143f308f43ef456041b;
mem[212] = 144'h010904c1f4650a8c0e11f611042e017ef507;
mem[213] = 144'h07d4f044026801790586072f064bf491f195;
mem[214] = 144'hf7b9f9a7fabc0d0df3d1078908bb001cf74b;
mem[215] = 144'hf28606b5fd720efd091e0f470054039bf5b2;
mem[216] = 144'h0ad6fd2e0df3f06b06a10adbfa6df96c0a99;
mem[217] = 144'hf6c9f89c0dea0b4e0127f9b5fe1ef7b0f705;
mem[218] = 144'hf848f4f7048f0d32f7b8048bf56df096fb5a;
mem[219] = 144'h0eee0de2f4ecf02ffb4b006dfbdf0c8cf3b8;
mem[220] = 144'h07f007ebff41001e09980addf4020a41f71a;
mem[221] = 144'hf6fd0075ffb1f79df5bdf2a70e03f95b0949;
mem[222] = 144'h0e7105b009f90b6605ad02b003ea09470704;
mem[223] = 144'hf955042df6f8f6b1f05ef49cf0cbfb810297;
mem[224] = 144'hfdfbfc23055c00200a1af772f8ecffee0d44;
mem[225] = 144'h049404ca07c503da0de4f7d90bfe04cf0a6a;
mem[226] = 144'h0d140df00ad30186f1710698f591fec4f734;
mem[227] = 144'hf045f038f32bf79b00f404a0fbf8f95909cc;
mem[228] = 144'hfdc50d2ef0c207d7029f0db80489f73003bb;
mem[229] = 144'hf724f63002c4fdf901cc0c80f47903b4f758;
mem[230] = 144'h0a310c26f493001efebbf8fbf5a505720d2c;
mem[231] = 144'h04f605540c67f4d6f6d7f32cf020f743fde6;
mem[232] = 144'h0276fee803ff0424f0c90b0a0e450184f06a;
mem[233] = 144'hf36605fafcbafa6404800ca60c6b065d00ba;
mem[234] = 144'h06d0f6b70113ff5bf5e202400b6302cbff4a;
mem[235] = 144'h0459066efadcf5d0f1e5089afaad04a2fad5;
mem[236] = 144'hf0f60527fba60a560c80fc6fffde0a6c069c;
mem[237] = 144'hfee7fd650bddf8f6f453fa8f05c20094f273;
mem[238] = 144'hf0b30bfe017b08d1f2def9a20fd0faebf5e5;
mem[239] = 144'hf81001ccf830f85a0c9c02c20303f426f83b;
mem[240] = 144'hf4a60fa0013707b500c705d809e1fe6cfa02;
mem[241] = 144'h0f60f07c044af33c09060243fa44073ef7d0;
mem[242] = 144'h035107a7073cfca4f7b3f13ff1fd0cf50297;
mem[243] = 144'hfd50f202f9350e5d0dde0f420b8ff030055f;
mem[244] = 144'hf01303640e1007cdf4ba02a7045ef3ef00e9;
mem[245] = 144'h0e5cfc24fd60f64bfe6e0c7c053c095d0fa2;
mem[246] = 144'h014df8bc08d7f61f00ac0b920d38efd8f11c;
mem[247] = 144'hfdc8fb95fbc608bff72706470e2b0ea40831;
mem[248] = 144'h003bf9d0f9f9f590eff7fe0902b0039bfa47;
mem[249] = 144'h097d0d05fc200b880baefb8b0b16fd33f717;
mem[250] = 144'hfea4f537f70c0381f51806b0fda4f08001f9;
mem[251] = 144'hf7040298f5caf2380810093e01d1ffb20162;
mem[252] = 144'hf289fa910440f718076200ab0d97fcf3f3c3;
mem[253] = 144'hf1c9f8e7fe1b0a3409bff7a8f2c409290bde;
mem[254] = 144'h0477f62cfc86f22203590dd6f9edf0c50bcf;
mem[255] = 144'hf042f27c00eff611ff64f26c067af6860aec;
mem[256] = 144'hff1ef1eef60900b20b6bf54efcdbf6760fdd;
mem[257] = 144'hf963f386f72afddb02e9fb4100f5f59ff924;
mem[258] = 144'hfbaaf813f37bfcbcf04803b8fd03fc5d0335;
mem[259] = 144'hfde50d49011ff4580335f316f7fd0dbcf8fd;
mem[260] = 144'h054407900641f8750425f07e0f97ff86f61e;
mem[261] = 144'hf058fde10a6ef67afa560930feb70a080993;
mem[262] = 144'hf64003010bf70397036b096cfa37ff880196;
mem[263] = 144'h0464f59ff42dffde0720f420fe3907c70d27;
mem[264] = 144'hf0a50b6501d6029df2670d8efd9b00e3f91a;
mem[265] = 144'h0030f2cd083100790ee1fa4b048ff4a6fa19;
mem[266] = 144'h0051fa0df989f9a407cef5870e58f175f5c9;
mem[267] = 144'hf81802890e7f06750fae038bf348f378fbd6;
mem[268] = 144'h0249ff1f042902f00d22f3abf691ff0ff8ab;
mem[269] = 144'h0933047b01cc0d46f9dff891f318fa8d0104;
mem[270] = 144'hfe87fc3df80cf715095c0cc4feec0bf106fb;
mem[271] = 144'hf8e10277fc840722f53bf7be00a40092fb0a;
mem[272] = 144'h0a07febbf42e06750634f7e10d68f0d3041a;
mem[273] = 144'h0b3df9a00eff00b8f965f0dd06db0fd8028f;
mem[274] = 144'h032506e1f522080b05570530fe95030ff80b;
mem[275] = 144'h08fb0cc8f027005e032af5c6f0b4034ff452;
mem[276] = 144'hf83006d101bcf369f5b2f964fc600bf8084f;
mem[277] = 144'h09bf0c5df4c9f2e1f2ce00e20d67fbc8f122;
mem[278] = 144'h0b55f85f0a600bcaf16dff29f8bd00d6054a;
mem[279] = 144'h0056fdeefd81071706c9fa180f6cfc3d000c;
mem[280] = 144'hf021018cf28d00e1f926f50ef671f098f39b;
mem[281] = 144'hfe0df962f4ef0d400245036b0ef00a04f6ab;
mem[282] = 144'hfa6a03dcfbb3085dfcfdf1700363fbf508a9;
mem[283] = 144'hf1d801690d46f5f0062f05ef0e8af41705f6;
mem[284] = 144'hfb2df1870c83f27ff7020a2f09e4febcfeb9;
mem[285] = 144'hff3ff128f0a408b7f635ffe9088d02a3f1ca;
mem[286] = 144'h0375016902c2f0bafeb901250a8807a2fc81;
mem[287] = 144'hfc3d01db0a1604ec0618f08c0dc606d5fa00;
mem[288] = 144'hf6a9f6fdf3bd074cfc3c03da0246fa08fa24;
mem[289] = 144'hf6bcf93706960aa40381f170f536f40ef1a5;
mem[290] = 144'h0564062af98000b70cf4f130f67c01e004e3;
mem[291] = 144'h0a7e0a87f8f6f153049af0380ff90c88f7c1;
mem[292] = 144'h02f10614f974f186f2a7f172f860048603ae;
mem[293] = 144'hf62a0dc4f362f025fa8efac80c3d09eb013a;
mem[294] = 144'hf6fa0d25fc26fd5ef0930f000670f9b60daa;
mem[295] = 144'hf41e09effc7a08fff741fd24f756f94dfbfd;
mem[296] = 144'h057101a1f7dafae40b61f036f5ee01100b1e;
mem[297] = 144'h029608a40b0af8e4086df61f0b90f313ff32;
mem[298] = 144'hfcb2f1e40a76faa1f7220fca041905b40239;
mem[299] = 144'hf1a9fe570de109a4f9f1fb37f32cf28a0e64;
mem[300] = 144'hfa1df7f7070ef130fcb30bb0fee8f3c5f328;
mem[301] = 144'h0c8bfaf1020c0e470c7dfc8ef00401e9f6c3;
mem[302] = 144'hf29cf7c6f01c0f7409dafe51fd0efc96fa53;
mem[303] = 144'h0c210d510f56099f041bf0640f1cfeedf7d6;
mem[304] = 144'hf04a052a045f0eeef1ea04500e7af6e5f50e;
mem[305] = 144'hff070649f274f27af2eaf0fbf4d505770c9c;
mem[306] = 144'h0c9b08b4fd8affaf024ff01b0bd30b11f1e3;
mem[307] = 144'h02d90d2802adf9ff0d790ad30361fd7505ed;
mem[308] = 144'hfb730d6ff15df8d5f6d8096efea6fe57f4dd;
mem[309] = 144'hf82003490083f5c10ae6f8d40696f1b9f847;
mem[310] = 144'h03380315f60d0d9ef36b00e20e440b260f63;
mem[311] = 144'hfdb4f4d20f700e67fc91f097fb860c970884;
mem[312] = 144'h0b2bf292fb0d06b3f2b20aa5f027f0560f1b;
mem[313] = 144'hf9fc008efa890d730677fa6bff200bb0ffe6;
mem[314] = 144'h006ef6760a54f7c606190bdd0b8700960fc8;
mem[315] = 144'hf01afe3efcce002ffad2f24bfbe40d130f94;
mem[316] = 144'hf79207b8fab50e31f4800ac9f73a074cfa24;
mem[317] = 144'h09790f1afa36f4f80e4df36b0a60f6d604fe;
mem[318] = 144'hf74403610b5c05e2f7060e62ff420f25fb45;
mem[319] = 144'h09d2f41dfa62fe400bb2076c0c700e57fb2b;
mem[320] = 144'hf9a30adaf54c083e07c0f615f62a0d9109c0;
mem[321] = 144'hf92df17407020239f82b083dffea0dcb0460;
mem[322] = 144'hf2c507b000e5f2d5f4edf48a02fbf9090e16;
mem[323] = 144'hf4530583f556fa49f6daff29f793fc90f20e;
mem[324] = 144'h01720f050b5204e400c206acf3a5f463fe8c;
mem[325] = 144'hfe29072a017404d5f29afef80474f2a9000c;
mem[326] = 144'hf794f4f5002e00bc017ef6850a35f1c0f545;
mem[327] = 144'h0f95f0700f24033e02a203c7f862fc56f5eb;
mem[328] = 144'h0b33fb2a0b8afb080cf5facc0adc0a4400c3;
mem[329] = 144'hf652039904070b730ee3f5790cd1003e0a6f;
mem[330] = 144'h012204b70256fc37fe2007c20d1e0daa0fa2;
mem[331] = 144'hf50b0728f7de07c20a51041fefec05f6080d;
mem[332] = 144'hf7a6f26c0af3fe57feb20387f2d800deff45;
mem[333] = 144'hf475f271ff570d6c00730cc9fa88089ef720;
mem[334] = 144'hfa04f88201cef4b606ddf3bffcd008eaf542;
mem[335] = 144'h0f60fda4f88900a30de6024300a2f2e9f55b;
mem[336] = 144'h095101d004b801c70ce10822f93908f70c38;
mem[337] = 144'hf45cfeb7fcfdf829fe67f105f207fd88fea3;
mem[338] = 144'h013bfa30f8cdf80600130b98f0ba0539f2f6;
mem[339] = 144'h02e308d2f5710e580c50fefbfde901a6fff5;
mem[340] = 144'h08fbfa860318040d05530127fb75f48405d3;
mem[341] = 144'h02830c8af53d030ff473f040f81509a7029d;
mem[342] = 144'h0cbc0d5cf8e30afc034df627fe6300fbf013;
mem[343] = 144'hfc2c09dbf9c7f9a6ffbeffe4f05cf05fff34;
mem[344] = 144'h081ffa9cf3270156f490f3e0f8e007f501a3;
mem[345] = 144'h0447f3b6f0eff9f90402fe9cfa4af51efb02;
mem[346] = 144'h0f1ff78ff04cf1e3049c0a1201a30e990e0c;
mem[347] = 144'h02a0f4fb0c32018bf6490a61f666013701b8;
mem[348] = 144'hf4d001e700740e85fc73fa230221076ef831;
mem[349] = 144'hfa77fbe00ea9fd4f003dfd100bd0fcec04be;
mem[350] = 144'h0867fc26ff230616fb7201f00c2ef8da07d8;
mem[351] = 144'h0d1600d903cb07d2f57400dbff570c010908;
mem[352] = 144'hf71f0853f24404b00e57031b0888fc2602e1;
mem[353] = 144'h068efe6b0e360c4bf82c01720cf8fcf1003e;
mem[354] = 144'hfdb500550a7efe52022af8d50cc80345faaf;
mem[355] = 144'h073c06310598f6a2f18f0d12078503130f8d;
mem[356] = 144'h01e2f308f097025ffeb002c709210f71f900;
mem[357] = 144'h02fcfb91f4ad0e1af90afd900683017ff172;
mem[358] = 144'h0460f35cf325084f0904f08ffcfaf031f3e8;
mem[359] = 144'h0ad2fb470dd10ca70e9ffb07f23cf4450298;
mem[360] = 144'hf7540ad9078cfee5058b01e1fcdaff060126;
mem[361] = 144'hff8901eb0428f3fe0177099e045f07ddf165;
mem[362] = 144'h0fb0f55ffdd002f10a270af70a3a0a1bf3a5;
mem[363] = 144'hf2b8f67bf71af03df8c0fe1c0ab10341f2f9;
mem[364] = 144'hf3fd0e9e093209ec08f70ff6ff72f884f5ec;
mem[365] = 144'hf23a0ba4f2adfa630ca00dd6f061f583f3a1;
mem[366] = 144'hfadafd3dfa0b05b300d9f5bf0cabf0d508b2;
mem[367] = 144'hfb8305fff316f549fb7dfc80f717f62cf288;
mem[368] = 144'h0a8a05cf0e4ef9f2f46cf1bef5a4f7eef60b;
mem[369] = 144'hff730085f534f611f7380fe40281f716fe29;
mem[370] = 144'h03bf08b9095e046af6060103fe7e050104d5;
mem[371] = 144'hfdb5f65d022affa809f9fd3a01da00330cef;
mem[372] = 144'hf9a609cf0ddcf669f6e5f6c0f9c30f1903fe;
mem[373] = 144'h0eeaf684f1d5047c0a7f06f907880ca20bff;
mem[374] = 144'hf49ff494f5f204c30e82faff0fa4052ff532;
mem[375] = 144'hf18cf7100995fb730c89f03ffc1a043a0b65;
mem[376] = 144'h00b7f9abf8ebf064f6cff6d006f0089dfa65;
mem[377] = 144'hf3470e9b08e0056901fafdef0df1fdc209bb;
mem[378] = 144'h09baf85b04caf8aa0cb10c52fe9bfd3afd9a;
mem[379] = 144'hf211f0aefe36f994fc5ef27a05edf6ad0e56;
mem[380] = 144'h01e80e30fd02fee2f31f02800655f8dd0440;
mem[381] = 144'hf280ff350df60234fe66fbdff7caf9bbf37b;
mem[382] = 144'hff47f6fbf1840f1e02f0f2fff6d60d45ff52;
mem[383] = 144'h08a5038e068bf465f1e6f49ffae8f968fc0f;
mem[384] = 144'hf78e0245fd29fe8b0dc3f247f098f9f1f798;
mem[385] = 144'hf86cfd17fdbaf1c8f06afdb5076c0e60f426;
mem[386] = 144'h01e2024df8c006b3fa5f00b6f1dbf9ea001b;
mem[387] = 144'hf6bffe790172fe3af109015ffe0902cd023e;
mem[388] = 144'hfebd05d8f050fd19f70cfd3e0761fdb90e22;
mem[389] = 144'hff2e00fbfda0fe5f01c0fd23085ef5f8ff56;
mem[390] = 144'hf7a90450f3ef0db9f63b0acbf9490150021a;
mem[391] = 144'hf5aa09f30dfff3ca0729060301ea01810570;
mem[392] = 144'h0057fa85f3b2f430fa5f04fa0b4c025c0181;
mem[393] = 144'hf2070745fe030913f66ef2a9fce9f50805c6;
mem[394] = 144'hf786f866f1acf4910c5805e40f09f289f6c6;
mem[395] = 144'h01370c47fbc6f3fa0334f2dd06ff0cba0535;
mem[396] = 144'h00d6fbc70b990a7ff678065af0a0047c0f6f;
mem[397] = 144'h0b3ef2bc08d8f0a6fc44fb36092b098b0bc4;
mem[398] = 144'h0c17ffab08a209b4f8f6f3b100d1042a0a87;
mem[399] = 144'h0cea05cff1930c31fea0ff8104ce08af0ac3;
mem[400] = 144'h07d3f92303d9f6b0f0bc0efc0d370c940123;
mem[401] = 144'h05650711f1560046f67cf8fcfa9102c908fa;
mem[402] = 144'hf7240e7403b00fc106c90225f334fa7b00ea;
mem[403] = 144'hf85f09040ec70a41fd3a0642034af40c0849;
mem[404] = 144'h0d76f58b0482f8f00c75007f04a308310223;
mem[405] = 144'h03dc0da3ff72fbd5fa040316fc9b0a7ff5f3;
mem[406] = 144'h08d0f814f788061efe9ff871f97dfdaf01c9;
mem[407] = 144'h0674f35003d1fb74f2b2faf7f750f7f9f62c;
mem[408] = 144'h03cc09820aa90611ffedfd05fde9f9eef598;
mem[409] = 144'h07030d81f358fc39055c025a0c4ff27d0a20;
mem[410] = 144'h0e0407a906c304b2fa3efce3f026effb0c5c;
mem[411] = 144'h0a33f83bfc3e03b3f8a9f351003001ad0aa7;
mem[412] = 144'h07e0f50005f0f6cf09b60f7406af0b6e0a91;
mem[413] = 144'hf9c70f31fcd4fdcd018e0395f6430cd2f9f7;
mem[414] = 144'h0420ffc8f0e7f2250ded0d59064cfda501d9;
mem[415] = 144'hf95d0a6702df048ff2be07d2f6f8f1b20c57;
mem[416] = 144'hf123f64ff59cf7dff063fa40efeb0b280c43;
mem[417] = 144'hf22806e10a01fa1c018afc96fc86f4e4f621;
mem[418] = 144'hf358f57df33f0dd401b1faa80ff3f605fc21;
mem[419] = 144'h0fc8f00f041cf08f0307f287f5ca085f07e5;
mem[420] = 144'h0c5bff64093c0ab0f9a60ad30adc01df062e;
mem[421] = 144'h03c0f6b7f02bf04808f302e8f1fef2010f67;
mem[422] = 144'h0bdef0510205f74e0d27050afde20917083e;
mem[423] = 144'hf988f81afbc5fdf8fa190f6d02e8fcb30ddf;
mem[424] = 144'h002603370874fcc9f020fd5906d3fba80113;
mem[425] = 144'hf7c1f1b4f2abfc62f5e001ba03be0ba5f43d;
mem[426] = 144'hf12bf3fc025b0d6bf67e0ebcf2fc0158012d;
mem[427] = 144'hfb58f61ff6230355f016fed1025000520f23;
mem[428] = 144'hf525f2e3ffc30e18f01401e70267ff750338;
mem[429] = 144'hf611fb22f187fbbcf6fbf81b06590b8f0f6b;
mem[430] = 144'hf215f826ffa40f54fd78f2c30a63f1010db2;
mem[431] = 144'h097a0041070c0fb1089a0a5e0308f261ff3c;
mem[432] = 144'hf6c3f94c03380ec3fc3102bafe6cfceb0378;
mem[433] = 144'h056af41ffac60c320ce80b4303bcf3f509ef;
mem[434] = 144'hf0430d070570f2f3f48dfd2f0bb5f334089a;
mem[435] = 144'hff4001b2fa5c093bf64b004c09c104b30639;
mem[436] = 144'h0c240e0f00d9083cf7f9051d00a808360f50;
mem[437] = 144'h03910f4af842f6eb0bf90f24064803020cd1;
mem[438] = 144'h01770b190737067cfd20f534fdd5f4eaf376;
mem[439] = 144'hfd6209abfcf50676f59d09ef0c63f5750303;
mem[440] = 144'hf9dcf30e086ff700f14b06960c34f531f76c;
mem[441] = 144'h0643070e03d70b1a0465f0faf2c408adf1a0;
mem[442] = 144'hfd7cfe91f3210d93f1b309530c7c0378f350;
mem[443] = 144'h007e0ab3f82c05c009880a81f9f1f37cf573;
mem[444] = 144'hf48209eb076cf9770c9efd120201f5c4f674;
mem[445] = 144'h0476fc93f5940d27f08bfd41f2970d800f2e;
mem[446] = 144'h026cfdd4ff27024ff70e03e6f4adf31efc59;
mem[447] = 144'hffa1f4b30ca7fa6ef115ff37fe55fa0bffca;
mem[448] = 144'hf8b1fd87029c0d5206b708d0fd440370f57d;
mem[449] = 144'hf76f03d3f0fb0d6905bf0934fd3908f50d49;
mem[450] = 144'hf1e3080ffb1d0e83fc2bfd4103a3f926f90a;
mem[451] = 144'h0a44fdcc00a4014e0975ff8109f9fb1e059a;
mem[452] = 144'h0f0df46bf9510bb40cacff64fc340f3a0cc5;
mem[453] = 144'hfbbcfd1afadefe2e0243f8c9fc6df1c503e8;
mem[454] = 144'h0c7df9bb0817f795f958f931ff19f4ba075b;
mem[455] = 144'h00def98406cf0c67f32afdc104c3085b04ca;
mem[456] = 144'hf0c107a2f2eff38a0c0a0d3203fefba0fe55;
mem[457] = 144'h0144f273f9d9fe2bfdd7f51a06ccf8570aa3;
mem[458] = 144'hfc9c02cd020cfa6e0b5105a70b780b5df816;
mem[459] = 144'h00d4f42e0e68f1dff00cf72efd460dc20d4b;
mem[460] = 144'hf331059bf2db0d650201f0500f9307eaf87d;
mem[461] = 144'h067f03d90d4ff8bffbaefac30a46099cfcd3;
mem[462] = 144'hfe4bf4240007fef2f6a8fdb7ffed0a73fb70;
mem[463] = 144'hf2c50cb5f65407aff6d1f06b069ef7e2035f;
mem[464] = 144'hf4faf476f0fbf2a2050609f9f601ff45fe34;
mem[465] = 144'hf6f0f32ffd50fc7cfb510afb0584f9bef80c;
mem[466] = 144'hfa50f926056cf535fcb00f7cf0dcfb5904c1;
mem[467] = 144'h0349f1b70b89f174f6bb0b45ff92f9fdf8f0;
mem[468] = 144'h0812051b041bfd54f3d00b4903d0f15704c0;
mem[469] = 144'h0601f87ef041facf01c9f13f0a8ff75dfbae;
mem[470] = 144'h0e2b0ce4f4890141f810fb9ff60209e200e2;
mem[471] = 144'h088406420428f36ff8df024c0017093cfbdb;
mem[472] = 144'hf143fae30690fda5f20904710f760b6df7a6;
mem[473] = 144'h0868070b0b080a6d05620d5bf3e8f8f5092a;
mem[474] = 144'h02f70ae7f4e00dcc0a3a0d95fce0fb580c6a;
mem[475] = 144'h0b29059dfba20d7ff63f06a30e4ff2a60aa1;
mem[476] = 144'h0df2fe86f45ef9c1f4b40f76f60d014e0191;
mem[477] = 144'hfdb500650417fbd1f19fff49fdc5fd1e0eb5;
mem[478] = 144'h0f920565007ef67cfb92f14400affeb1f338;
mem[479] = 144'hfdda0e9c046d0e71fdd6f78406c5f127fbc2;
mem[480] = 144'h0704ffe80f58f2c60194f8b3f7880b1a0a92;
mem[481] = 144'h0eb70a6af8def8bdf847f5cf0d1107100dd1;
mem[482] = 144'h08e3040ff9710f0d0268f1c1fa1e01110d80;
mem[483] = 144'h0a22fe030fc6006df568039d07ecf8ba029b;
mem[484] = 144'hf07ef635fd9d07c00532ff2c0358fb3b0f74;
mem[485] = 144'hf98707250664f47b06bd0bdbf7aaf6fb0daf;
mem[486] = 144'hf96ffe8df3d1fc100a9e04e6ffab0f72fee0;
mem[487] = 144'hf760057d021f0bdb0fbd0f14049dff40fa66;
mem[488] = 144'hffc0f862fe9cf98f0303fa8ef594f1660b5b;
mem[489] = 144'h072ef14ef2880ab80ae0fc3c0b1703640f9d;
mem[490] = 144'h0e1e0bb7fe8bfd70f375fd78fa220aedf843;
mem[491] = 144'h09f30ed7f008048f010c04080deef5c8f916;
mem[492] = 144'hf040022905f2081e070c0219fc21fe0af136;
mem[493] = 144'h0bc9fc90fbd80d2b096c0183f9e2f9ecf391;
mem[494] = 144'hf434012bf9980af107d40f11fddd0638f3ce;
mem[495] = 144'h0207005bf15608adf4c40d8ef22109a10787;
mem[496] = 144'h0065014c02a10483087d066b0307090a0ab8;
mem[497] = 144'h0ce50ba60eacf9240b5600540c5ef39ffc4e;
mem[498] = 144'hfaaffeca05c2031af09efcb0fed60fb4fa93;
mem[499] = 144'h0e7e0ad90acafe4203a3f3befccaf4c203ca;
mem[500] = 144'h0fc1040c017bf239fa73f8b20123ff40f53d;
mem[501] = 144'hfbed00f30b1ff2d4faa00c650e92f8320cb9;
mem[502] = 144'hffdbfa71f5310440063602130be1f91502ee;
mem[503] = 144'h0403f8ef09ecf2c2fe0c0de80848f299f0e3;
mem[504] = 144'hf1a3f774f2eb0472fae106f5040d0eacf188;
mem[505] = 144'h01c3029a08370c8e094e0092f16ff172f0d6;
mem[506] = 144'h019606f1073302d80ed3ffbdf76bfe750b2d;
mem[507] = 144'hf208f0bb0f3d095df696072100b303630034;
mem[508] = 144'hf67b0d1706f8fb0c06cefa08045ef2bd0ef8;
mem[509] = 144'h0c8d0eebfa17f24f09baf9c30abffaf3fa22;
mem[510] = 144'h05d20264fe9503570e70049203570a01f827;
mem[511] = 144'h022605b80fb704aff8ebf8bffeb9f3c20e08;
mem[512] = 144'h0d9afa4d041409d1f63f016402bbfc2805f0;
mem[513] = 144'h0f760e0eff9cf539f42dff1ff453f429faf1;
mem[514] = 144'h03c3f3f5fc90f7a70261091ef329f0e50a00;
mem[515] = 144'h049203b1fb08ffb30df20365072cfa7609ee;
mem[516] = 144'hfe9103dcf61b0ea8fa6c0750075cf5990050;
mem[517] = 144'h0830fbd1fd49efe20dc5fbde0cd702eaf193;
mem[518] = 144'hfc3d0f85fdcd0f6df0080059f5a204a80f55;
mem[519] = 144'h06ccf63af4a3f6abf64200fafa5103a5fdcb;
mem[520] = 144'h0ba40b0702a5f27f0d1df6a305b6f04df5ed;
mem[521] = 144'hf891f96e05f807d00846fa24fb680a7a081c;
mem[522] = 144'hf8170af0fae2f6e50971fe3df79a082ef743;
mem[523] = 144'hf7340117f37a01800ebff6bf078cf2bc058d;
mem[524] = 144'h04670ce70bacf6eef233074af40402bbf67b;
mem[525] = 144'hf48bf833f03af32401820f5efe30ff920fd2;
mem[526] = 144'h0a3bf78ffe0ffa6900b5032c00d0f95bfa12;
mem[527] = 144'h0f340b98f169ff94ffe2062dfb1c0a510c0b;
mem[528] = 144'hfff60d75f8a40cb6ff65f600fbbdfa7f0b6c;
mem[529] = 144'h0afbf38ff1770137fa0b095a07b60fb0fb9f;
mem[530] = 144'h0fc00191fc88f23f0dd102fd021506a40933;
mem[531] = 144'h03ee07b707f9051c0521f52af4b10a97f080;
mem[532] = 144'h00a7fe1c07d205fb0a660f04fc0afb630413;
mem[533] = 144'h0020fc2809f10985f3c1f4bffa310631f2ce;
mem[534] = 144'h0e4d0a00f97d08db045df1e2f01a09c7fbac;
mem[535] = 144'hf6d6f86af852f03a07b40d5d01890f140a3d;
mem[536] = 144'hfaab020e0a40f29e0539fa27f557ff990c99;
mem[537] = 144'hfb0cfd3d06830593018a010b0bed0ef9f542;
mem[538] = 144'h04e5f463f9810f6df278f0410e690a59070d;
mem[539] = 144'hfe39049af99afc23002bfae5fd6ef623f7e5;
mem[540] = 144'hfd63f3c1fa5af01100d0f626079f059aff01;
mem[541] = 144'hfa89f5f80a040542ff9b01a9f2910b06052c;
mem[542] = 144'hfc0fff4b05910676f6df06e8f186f9c8fdf8;
mem[543] = 144'hf594f82103180a8b03ecfd48ff1905f3faac;
mem[544] = 144'h0b60f7a6fa58fdf8f531f6af01ee0a010405;
mem[545] = 144'h01d8fa8b00bc0761f71d036ef821f56bfbdf;
mem[546] = 144'h04b90f01f69ff999f36bf9e7fa6c0cf6f3fa;
mem[547] = 144'h04920dd20dfd002bf6defc93002ff752f6bd;
mem[548] = 144'hf2d80516f6cff84d019bfc05f3e50c6e0999;
mem[549] = 144'h0378f6be0f79f9410935f52f085b0d58f768;
mem[550] = 144'h0de0f93a012806b909da08a9f6bb0a06f899;
mem[551] = 144'hff7ff4e4fbcdfc6f0f0408220825ffd304b6;
mem[552] = 144'hfd5bf742f47c0975f889f50ff48bfc0c08ab;
mem[553] = 144'h083d0e77f4f9f3a7f0240597005407d0f99b;
mem[554] = 144'h012df429f1370f5d06690e0a03a3ff72f4ea;
mem[555] = 144'hf458078df1470af7f17e03b30e00f19d0665;
mem[556] = 144'h0e84f2e8fff90fd4f5edf92e08f8089c06ae;
mem[557] = 144'h0039f3a6003f04e605ae0387f33cf311fd19;
mem[558] = 144'h035ef4d0f9ba03defab40e7c02440261f773;
mem[559] = 144'hf59007ddf95b02ad089df8ee0e91fc91fce6;
mem[560] = 144'h05f3f9a5ff3808a10cc9f610f1e7fc3efbba;
mem[561] = 144'h0f47f25a0ca90767f7070b29fbb50695008c;
mem[562] = 144'h0145fe26072f0a08076d0cdbfe6a0bb4f509;
mem[563] = 144'hf1fcfa68056007bd0d3c01090560f2370f9c;
mem[564] = 144'h091ffe4ff334078a04a2f7a2fbbdf236fd5e;
mem[565] = 144'hfcdd0b0bfddc06c3fa8ef535082c04fafab3;
mem[566] = 144'h07790c080d940af60529f0f6015ef9c3fa7f;
mem[567] = 144'h0c59f858f34c059100240f51f4d8ff390fd2;
mem[568] = 144'hf017f8ba0bbd07b1fc98f628f48d05f8f44b;
mem[569] = 144'h01eef659fa7cf0f109e5fa9902c80d93fba5;
mem[570] = 144'h0859f86e0153f7c3099a090bf1d40210f253;
mem[571] = 144'hfe0602d702660eff0e3dfe0a06aa0b51f41b;
mem[572] = 144'hf915f8ce054cfd4ff65efa6df05b0a5cfcd6;
mem[573] = 144'h0c9a041805340a770ed2f0a20f6c0207f6c2;
mem[574] = 144'hf05cf3d4f60ef7bcf90b0ba6f244070b0b63;
mem[575] = 144'hf5010ef7f057f8e6f639f8be07bd03b8f5ea;
mem[576] = 144'hf70508ee089f018df8dafd71f09f0940f916;
mem[577] = 144'h0cd5fe5e0f9a0a030b420906010103b90675;
mem[578] = 144'hf76b02e90a37f2740f0ef2fa027df3d0fd47;
mem[579] = 144'h0dd707a8ff4a0e34fc2a0c00f4e1ff9a0a0a;
mem[580] = 144'h06f70b400cafff500b0bf7c209f1f2f7f1c1;
mem[581] = 144'hf651f2120e93fdfcf37002d202e5040c0b1d;
mem[582] = 144'hfafff9eaf7e4f82ffa7e058e00b9f2240c37;
mem[583] = 144'h0fe0f3aa0776090a0e6efd2e0d110fc602fe;
mem[584] = 144'hfcea0c570edafc22f4cb0b2af2bc019bfb3b;
mem[585] = 144'hf388ff9507db036709d4f65b0639f332fd6c;
mem[586] = 144'h0590f808f6fc085efa040ebc067cf7d30276;
mem[587] = 144'h0e050cb4fb4af244f98dff3c00e709aef22e;
mem[588] = 144'h0c2d0096f2bb04d5062f05c609c9ffd5f820;
mem[589] = 144'hefdd0ea60f7bf4b6057e0d050370f7e00e81;
mem[590] = 144'hf9450915f54a02e9f00afb370174f128f972;
mem[591] = 144'hf98905f6090c09560b730dbcf22f0773fd87;
mem[592] = 144'h0637f3e70b160717f20afd25f0ce01a40ce4;
mem[593] = 144'hf37604b7f56df59af34cf67805010416f91d;
mem[594] = 144'h0786f35a0d99fb55037bfa35f2380e9005fe;
mem[595] = 144'h0c9f0bebf91b0994f11a04fbf1f0f3ed0437;
mem[596] = 144'h017306a20a500be20306f09b0cb9f695009c;
mem[597] = 144'h0022fb9dfdcbf93f015b0b36f494fcc6f074;
mem[598] = 144'hfb250ed10315febc0e960c84088c03bc08d6;
mem[599] = 144'h091e0167fa6400850d5af5b6075f06e7006c;
mem[600] = 144'h063b006af2db0f6607c6f58f0d420c6a014d;
mem[601] = 144'h030bf2dbf39c073504a0053f0ba10ced0d2d;
mem[602] = 144'h003af4140ed7f14903f8006bf84a0d6efad4;
mem[603] = 144'hf97e0d9c03e30538ff81f82f0fd808c70136;
mem[604] = 144'hf1e3fb0a0878076efa1708740e46fa0ff848;
mem[605] = 144'h0e8401c60d5906ba047f03f1f913f3f300bd;
mem[606] = 144'h0864fcb1f0250cb8fca3fb460197f77bf6bc;
mem[607] = 144'hfa430900fc87f530f07af9e6006706cdfa77;
mem[608] = 144'h00cb02090daefbb2039bfa08f2c0015e0727;
mem[609] = 144'h006ff0ddff40fb9306f2f7f4fb6bf0a30bb5;
mem[610] = 144'h0c62f660006af43906e20c2cf1d3fe170504;
mem[611] = 144'h061dfdcc02dbfe00f7300932faaffcdc05c6;
mem[612] = 144'h07cffdb60c3ffa4afa930f6afb1803aff44e;
mem[613] = 144'hfecef344f684f86004c7f134f143fb6cf837;
mem[614] = 144'h08eb0d87f780fb780113fbc90448f46ef733;
mem[615] = 144'hf4f904e302d101aa006a0c3f0ce9feccf21b;
mem[616] = 144'hfd6e0991fc380351f110f6a10b3b0204f447;
mem[617] = 144'hfd170aab0ba00e6ef18b0dfff67a0a39083c;
mem[618] = 144'hfd9d0ba0f17b0271f3840b47f457fee00deb;
mem[619] = 144'hf2eb03d30647fdc801f40d80f6e8fee705a1;
mem[620] = 144'h0afb03cc09c4077e0b85044cfece07a3fa0d;
mem[621] = 144'hf9def99cf64ff394fd6dfd5cf1c5f3360dc6;
mem[622] = 144'h0535ffd00eae074f0d0e02010c21002f0c06;
mem[623] = 144'h0ac2066af10bfc1df199f2e1f8f9f5b20249;
mem[624] = 144'h06930c4707c70ee5fbb7fd78036200bef65a;
mem[625] = 144'h020707f204bf0ccc0f58082000aa0c410a3c;
mem[626] = 144'h0b81f519f61af50ff9ac0506f9a10c0605be;
mem[627] = 144'hf9ee00b2faa2f2e30d05f3d9fe45f2e909ce;
mem[628] = 144'h05fe03d8f2d101d6f6c309aff082f8bffbbe;
mem[629] = 144'hf4440d21f657f8ce039c02b10b6bfe760707;
mem[630] = 144'h0973ffddfaac03b001f8039f05d109f604ad;
mem[631] = 144'h040efe0a0c7affcbfb450f27037bf06d0506;
mem[632] = 144'hf7010cc4086dfb790f280807fb6e067c01cb;
mem[633] = 144'hfd850479018b040afe30f41bfc310494051a;
mem[634] = 144'h0b09029e0066066df2a3049504b3049cf148;
mem[635] = 144'hf1210cda0c3803df0ca70895fa84062e0643;
mem[636] = 144'hf8d90bf4ff47f8970250f32f0769f3180ed0;
mem[637] = 144'hfb310c81fa860bd80515f2b5fcb00630fdfa;
mem[638] = 144'h0fa6fa3df3cc0440f5bb0b11f174f7b2fdf3;
mem[639] = 144'hf8440cfdf3d2f00cf32cf358fd5df30b06f5;
mem[640] = 144'hf6000b7a0b4eff7d0ad1087bf770fc7bf651;
mem[641] = 144'h04f9f9b2f4dc0d58fd570967f9cff278fb8e;
mem[642] = 144'h0318f1260346f1fdfea405ac00820b87f049;
mem[643] = 144'hfacb04bf0eb10dde0bcc00a507ff06d6f8e1;
mem[644] = 144'h038d04840667f7cc03e901f1f0ea07ed064a;
mem[645] = 144'hfeb8f10b082cf25a080df7ca02b80ad0f2bc;
mem[646] = 144'hfaebffa50536f9dcf3a205df06510f3ef0e8;
mem[647] = 144'hfa44ff6bf8fa0dc4044c0b4f04010058fd0c;
mem[648] = 144'h0bd90626f956085000090b07f2de0026fd72;
mem[649] = 144'hf3bff00a0bcffef0f987f99409620ff20ad2;
mem[650] = 144'h07a20e11f01900f4f6aef50dfec50d870c60;
mem[651] = 144'h020b0628f53b02be0645f9ef02aff819f2db;
mem[652] = 144'h0218f020fb54f48cf621054ff97ff68602ad;
mem[653] = 144'h01e7fa0dfa6b01f20d4cf8c9f5800c0df2a7;
mem[654] = 144'hff8dfbfbf9f3f66500a1f51f0099fd6e0261;
mem[655] = 144'h0dcaf7adf1c0fe75072cfa170cbc09910ca9;
mem[656] = 144'h0231f604006ef4f808520a4508c10978f48e;
mem[657] = 144'hfb02fcffffbd074c04a40e0304520c08049e;
mem[658] = 144'h04e3f884f6560674f17bff2a01fafb5df40f;
mem[659] = 144'hf26efed3fdedfc1b02840c90f42dfad5050e;
mem[660] = 144'hf2a20c68f572f42af86afc710b30f9c8f425;
mem[661] = 144'hff2af71c0dfd092ef508f6c2f262fc620b5c;
mem[662] = 144'hfa890f74f1970403000c08e2ff4b0c8c0ef4;
mem[663] = 144'h02f80e47079c0c5bf897f154fb370615f836;
mem[664] = 144'h0b10ff850bd706c80520fa2ffa68047ffbe7;
mem[665] = 144'hfab00e740efeff61fdaf0791ffcaf6c2f1c4;
mem[666] = 144'h00baffd808a7ffa1f4b201cff7abfb21fa90;
mem[667] = 144'h0ec6f073f055f46c0360ffc908b4062ffa93;
mem[668] = 144'h04a50ed30dfaf7ce0450faa5f19e0d8bf598;
mem[669] = 144'hfac8ff36080404e50251f7cdfc560f29f747;
mem[670] = 144'h0f8ffc88f74ff2e0fabe041ef3420fa30db7;
mem[671] = 144'h0f44fd060b340f790734fe96051d00f9f793;
mem[672] = 144'hffd105e40507f7740ba3fc080295f63ffca3;
mem[673] = 144'h0c2708acf877f8a90e760794f012f409fc08;
mem[674] = 144'h0d47f75dfd21f2c4fc54f485f7ba04320871;
mem[675] = 144'h00a2f5dd0ec8084901f1f37d0cd9021ff0f0;
mem[676] = 144'hfc100fcb0aa8f79a0f3804e10e10087e0925;
mem[677] = 144'hf159fb3d0b89f99d08bc074ff7e80c78f555;
mem[678] = 144'hfcf9fca20fa708ee0a14043cf916f5d9f3ac;
mem[679] = 144'h07f4f654ff4002acfadcf67a0c56f264086f;
mem[680] = 144'hfa47fd28f4e40094014bfe18f228f6380269;
mem[681] = 144'hfba0f72a03cb0bb80fdb031ff32c0fb4f036;
mem[682] = 144'hf40906cff4f8f7a90c1b0e410e51fb660f90;
mem[683] = 144'h0699f5870fa10766f0f609210c0f0c0d0a1f;
mem[684] = 144'h0bfd0b03f6af018ffcc709680c2c00a9f183;
mem[685] = 144'h009cf2d9f64bfdf7f48ef63afc9a0e090842;
mem[686] = 144'hf5e90749fb210264f767fca10eb40e5ef55c;
mem[687] = 144'hfd69fd80fac0f41708800129f319f476000a;
mem[688] = 144'h0b8df49af6c0f76c02a6f46ef78df271f2a3;
mem[689] = 144'h0d840d4d02850388f65e0284f89706effe8c;
mem[690] = 144'hfdd2fb520b4903bbfb830e5a0d320ba50aed;
mem[691] = 144'h0366f6fd056b09b6efd50411f6d804b70142;
mem[692] = 144'hfce7074d074cfb88f5220f900867f817f19c;
mem[693] = 144'hf2b10c43fccaf19b08aef5d40adf09b8fe3b;
mem[694] = 144'h01970dfc0cb40c40040005c9f3580d30f462;
mem[695] = 144'h0b5d0a8dfd09003f098f0a92f86ff2770bf6;
mem[696] = 144'hfbf3ff850e2ff35dfdfd0969f2bcfefc0b35;
mem[697] = 144'h0319f71bf8950a140ea2f193fc6af07bf1ea;
mem[698] = 144'hf376f1f40d4efc26fc630f4afef80838f805;
mem[699] = 144'h0d63fdfe0de0fc0e01acf492fa7c04090343;
mem[700] = 144'hff5ef2d3f2f70e33f03dfbf50384f7bbfa47;
mem[701] = 144'hfa6a0b05f9cc007df6ddf416f5c2ffccfdbd;
mem[702] = 144'h09bcfef8f713f9d60720fd3b0adb06ab0d4f;
mem[703] = 144'hf207f5670708f69206bcfdf9f146f80efdce;
mem[704] = 144'h0d470258f78506dafd47f0a00f5606ef06eb;
mem[705] = 144'hf096fcdf0ce40ddefb8afb30fa8df0770407;
mem[706] = 144'hf941f447fdb9f58ff9300c340a4ff09707e6;
mem[707] = 144'h0715fd03069309bcf40ef273fbeb04b500d2;
mem[708] = 144'h05ff002f08d405fe095406d70ee705780a19;
mem[709] = 144'hf9f6ff440e68fac00b50f334f2190a18f8e6;
mem[710] = 144'h0619f2b2095905aef3f7095e00c9f41806d3;
mem[711] = 144'hf1c1f95b0a46fb02f767fa23f32903cd015c;
mem[712] = 144'hf75401f3015ef360fc8b0da206e7f3020aec;
mem[713] = 144'h055308aef02e034103c503620c81fc6ff256;
mem[714] = 144'hfd9cf151fbf4f6df05c5fcf6fe40f416f111;
mem[715] = 144'hfccff113fb7afa3d00e0029f07b0fd0cf64e;
mem[716] = 144'hf5ca0c3901f0fce7fb2ef8a4efedfd56fab8;
mem[717] = 144'hf51c02def4b505690333044ffb2a0242032e;
mem[718] = 144'hf6c304a509f70c1afbb20a310555feddf540;
mem[719] = 144'h089cf38afb13fd17f0fd0c570aad0a9a0f3d;
mem[720] = 144'hf46c0018046505adf3c508840a70f2a4049d;
mem[721] = 144'hf247f15409810868fb83f259f2f0f32d034b;
mem[722] = 144'h04360fd60d9504d80a22fdfffe39f2750e39;
mem[723] = 144'heffef0810e8c0310f6defd27fd8a06710bee;
mem[724] = 144'hfcf5f190086ef13f0d94f346ffc4f4380bbd;
mem[725] = 144'h0fdcf6b6feda0b5f0127fe820a030b830186;
mem[726] = 144'h0aa8fc47f287f6da0113fc2401bdf175fa7c;
mem[727] = 144'h036f049300c8f55ff5e80c40fa4dfd18fe3b;
mem[728] = 144'h0df70a5a0abaf668f720fe06fd2a0e4e0910;
mem[729] = 144'hf6e90fb00e740204fb2df7edf4de01d90c94;
mem[730] = 144'hfe8a0da2ff8a025904f90e6408f101d60bca;
mem[731] = 144'hf2c4f48d07e9f071092cf87ef375febf0dca;
mem[732] = 144'hfb28004af549f2d8fc080bfd0ed5fcd8fea4;
mem[733] = 144'hfe7d06ec04a3fb87f42bf5b4f994003f0144;
mem[734] = 144'h07df0377fc3bff600df40db2fad509940e04;
mem[735] = 144'hfc750abcf3b20a4a07860ed0ff9bf4c204ea;
mem[736] = 144'h0beff387030ef3e8f401fce5f41305010823;
mem[737] = 144'hff6b04b8fb0bf99cf5d7fa3d0e7b0a17f303;
mem[738] = 144'hf96f006dfbf0fff5fe6a0ab30f6dfc0e0d6e;
mem[739] = 144'hf55807e80e11fa660a6406a70f0af96bf5f8;
mem[740] = 144'h01bef376f1d30607feebfe5001c20e28f64c;
mem[741] = 144'h039ff9f2068af4dc02fdf6140c37fa9c0ef5;
mem[742] = 144'hfeb707260da0f6390e3df1520a17054c059b;
mem[743] = 144'hfd11ff54ff0d048a0bc4f41300bafd5a0dc8;
mem[744] = 144'hf51000460a810673fa40f4ec0077fb9af4b6;
mem[745] = 144'hf49d0144061100160de5fb40084601d4f964;
mem[746] = 144'h0adff02b0cc60f43f8e402d9ff6ffbe2035c;
mem[747] = 144'hf70c060df094030df5fbf2c40e36f077f50a;
mem[748] = 144'hfdd20d7207a4f8cd07150f630492f6f001b4;
mem[749] = 144'hf7b1f7dcf6fe06580781f472f2f80e3c0702;
mem[750] = 144'heff906cf08e6faa209cf069df1e8f0daf77f;
mem[751] = 144'hf19406a8ffa20db6f422f8a00e31f641fed4;
mem[752] = 144'h0841ff250cf2fa550d00fd86fb51fcb4f644;
mem[753] = 144'hf29bf30e075b0129f7b602070c9502eefe15;
mem[754] = 144'h03e7fc690658f91a09cffa670281f4c6f723;
mem[755] = 144'hfed2f1fc0aae07f2fc67f336f5a9f2bc0dce;
mem[756] = 144'h03c80b770383f85803a2062b04dffe3a036f;
mem[757] = 144'h082e0cc6ffb3f9e7f86bfbe7fbd5f206f4c2;
mem[758] = 144'hf5c807e001ccfd23f27ef347061ff416f341;
mem[759] = 144'hfd40f1f50b8bf4d3f0570e85f5ca0148f2ab;
mem[760] = 144'h0414f68dfc85060404990992f8a40b6b03b7;
mem[761] = 144'hf3f0f348f4d80baef46df0bb0f49ff05f3bd;
mem[762] = 144'h0cdffc72f80bf46a0a7cfaf9f3dffe5eff5e;
mem[763] = 144'h0b3c03030bdffab4001800b6f724f1e5fa9d;
mem[764] = 144'h0359f64e0e8ffabbf15e0eddffa4045d0ba7;
mem[765] = 144'h095d019af7acf7180050ff5501e5f139013d;
mem[766] = 144'hf7fd0b1dfbedfc9af04f03ebff9501c5ffd7;
mem[767] = 144'h0139f32b0711f93e091a07ebf37d02660b9a;
mem[768] = 144'hf69004a80d55ff06f380fb2af052f8faf876;
mem[769] = 144'h0a79fdcffbb3018c003102eb0e60f8320964;
mem[770] = 144'hf185f7fe02d60a930949fbc3f780f1170050;
mem[771] = 144'hfb94fdd0f4f7ff3ffa2d09eb0c3b04450f3e;
mem[772] = 144'hfd5b0d4f0cc00b69fd22faa70f23fb740fe4;
mem[773] = 144'hf8d5f039fbb300fcffddf5e1099cf88a0bc9;
mem[774] = 144'h0f18f584f959088bfdf9014206a0f6fe01e9;
mem[775] = 144'hfbefff76f42ef43c0a01f764014ff264fbc6;
mem[776] = 144'hf477ff9df86a0b200735f75c07270f54f5a1;
mem[777] = 144'hf83af1cc044d0582f8bd02b2f501fe31f4c6;
mem[778] = 144'h047efefa0304f37a0bf70f2309c9feeefc98;
mem[779] = 144'h034dfffa078cf7dc08450612f818f354f002;
mem[780] = 144'h02780704f72f020a0d460712f5b7f8d6f749;
mem[781] = 144'h0ea4fb44f5290d4efbeef1e8f5b0f5b20854;
mem[782] = 144'hfda5f3fafd6504eb0b6102fef73a0ba70b33;
mem[783] = 144'h0097ff9df606f901ff9cf6bc02c20917ff60;
mem[784] = 144'hf00bf9eefea7f660f64a0c96036100fcf20e;
mem[785] = 144'h0ea0fc73015804ed0762f2f9f5b7f0850980;
mem[786] = 144'h0fd3fbacf33a0a30f90d096f09f009080935;
mem[787] = 144'h0e77015e0a92007ff8600468019ef886fa99;
mem[788] = 144'h0b09057e008401790f030d7e0cebf56ff15b;
mem[789] = 144'h00fdf58e03a401420fb80c6009eaf2f6ffa1;
mem[790] = 144'hf814fb93f059092c08fd0b0bf5db0515f3eb;
mem[791] = 144'hf7c20459f3f4f352fedef1baf960023ff10f;
mem[792] = 144'hf4fff11008b603c2f0c8f0f30bcbf9d4fed4;
mem[793] = 144'hf0fff73cf68af93cf898f2ce0cf8f673084f;
mem[794] = 144'h08e8f91c0a27032ff940fe76f604f5c10eba;
mem[795] = 144'hf185079205fe0b71f1af01f9071c05d30e74;
mem[796] = 144'h00340596f92803be0dbb020bfc7206530145;
mem[797] = 144'hff3a0e670f4d081ff18d0833f45104ea0ebe;
mem[798] = 144'h09fd0f2706a9f85c019d045d0e20fd00fa19;
mem[799] = 144'hf6820fe9f925fd20f5520032f848034c0fd8;
mem[800] = 144'h0e48fa14fef20705ffc501740b390cb5014e;
mem[801] = 144'h0e610dd301f6f95afde20385f7b00bc8f844;
mem[802] = 144'hf699fcc4fd320e05f22ff32bfe3dfa7300b7;
mem[803] = 144'h0d9a0362fed0ff5cf97c0c83fa0f0c6e03db;
mem[804] = 144'h01a5fecb0032feba04e10434f0cdfff8f471;
mem[805] = 144'hf07e086104ca0964f423f69af57b054202b1;
mem[806] = 144'hfeaa04f3fd39031af50500cdfa06fa17f7cd;
mem[807] = 144'h0003fc18f3ff0a08fc7302c60eab0a5ef13f;
mem[808] = 144'h0b5cf0c90a8a0906fb10076ff56d0a9df140;
mem[809] = 144'h0af9f9ad0db90cc105320536fb1ef60cfccb;
mem[810] = 144'hf60b0b1bf39bfeecfcddf921fdd6fb0ef0fb;
mem[811] = 144'h0763f97102cf072cf8da008308e5085eff91;
mem[812] = 144'hf7bd0598f7ce0c6f01a70112034ef9b800bc;
mem[813] = 144'hf562f33506c9f0930e9ffeeff64cf5dd021b;
mem[814] = 144'h0a96f6780f720e92f25af5b504fd0714f180;
mem[815] = 144'hf19af61e0b7f0a020e71ff52fc58f4b106b4;
mem[816] = 144'h0805f49df579f0ae0f2afdb4fba107730100;
mem[817] = 144'h063107220e98fbe3fc7c0abd042df78309cb;
mem[818] = 144'h036f0da40d97f002f1c10e74f7ff0a2803c1;
mem[819] = 144'h0ea8fdf5f98efd91fdb303e50ccbf99b00dd;
mem[820] = 144'h0a050ec3f82ef4e208af0dd40260fe78f722;
mem[821] = 144'h0a5af59ef6d8f1f1fa94015e06370e3cf01b;
mem[822] = 144'hf12104160ffbf51f062b0d13f52d0014023e;
mem[823] = 144'h0f4cf86204e3f36cfd4b0cfbfb3bf97b047f;
mem[824] = 144'hf65102e2f89e0413fbe2fa79fcaaf1790b00;
mem[825] = 144'h074709fdf747f1e7f253023f061f0b450416;
mem[826] = 144'h05e0fe9801240d080a09fc96003c0aa3fc17;
mem[827] = 144'h027cfb07053ffc2bfe4df9d7f1f3f6390f4c;
mem[828] = 144'h0114f130ff76f58bfdb100bf04dd08e7f5ca;
mem[829] = 144'h0641f3d5fc76fc1bf1690617f05df2d3fc9a;
mem[830] = 144'hf466f18a05d4094d07090f50fc55f06203b2;
mem[831] = 144'hf89002a80a6eff7e023501430e73f8f3fa92;
mem[832] = 144'h0cd509e2f59df79df8cffcbc0e8a0c40f945;
mem[833] = 144'h07b0057ef4340963f9b7fddc024a0f080e99;
mem[834] = 144'hfb1fffdaf1c7047e0466f00c0e92f58e01dd;
mem[835] = 144'hf69bf29600bcf5a1f628fd43015406e0feae;
mem[836] = 144'hfa17f28e0f17f82ffd49fda10757f21e02a8;
mem[837] = 144'hf79c003601d90af7f07bf547052004fdff7e;
mem[838] = 144'hf43507290577f600fde2f2cf07ae0113f02d;
mem[839] = 144'hfe9d03650f4bfb88f9c40a84fddc04990050;
mem[840] = 144'h0ea9f69207e0f3b3f3bff2effcd90bc70118;
mem[841] = 144'hfd200b5ef4ce00e9f5580d6df24d061bf26d;
mem[842] = 144'h06c3f6770a420608f1990f720001f06b066b;
mem[843] = 144'hfc7b05f50170fecd0628ff3b0ef1f1a70173;
mem[844] = 144'h08bb09e6f67809b30d49fcd40b4d0a35f5f6;
mem[845] = 144'hf9f50020f28207cc0e07f94a0b54fe3af344;
mem[846] = 144'hf9d00c350b6df332039efe83f733f8780258;
mem[847] = 144'h0d66fcfa0ca6ff150fa0f4ef0746f847054d;
mem[848] = 144'hf091fbf10a95f1ac0877fc9bfc130529008c;
mem[849] = 144'hf9aef46305c8ffb9fe0e011409cc00b80c61;
mem[850] = 144'h06f70378fc4af03cfd91f972f49005a20764;
mem[851] = 144'hf519f9020a8bf8fa0212048ffec4fa7dfb5f;
mem[852] = 144'h0b7ffc590298fc88f4c5f99df4da0c690579;
mem[853] = 144'h04ccf9480e6a0dcb09eefe3d0f98fd1e0734;
mem[854] = 144'hf265054c01680b610a030b6c01ecfe75fec9;
mem[855] = 144'h0f13fd3902d2081cff3f0d940b04f45601dc;
mem[856] = 144'hfb77034c039bf735f564f7500089fa950d5b;
mem[857] = 144'hf490f4730f5f002d00acf898fb4cfbe90676;
mem[858] = 144'h08330aa90487f084f2fef3b903d904ccf6b7;
mem[859] = 144'h0b71f0fa023bf3f5f36d0aec009e01f204c2;
mem[860] = 144'h017ffaa0fa71f24f0f4ff4feff4ffcd20fc4;
mem[861] = 144'hfaa5fbb0f45a006ef505f3a20348f98d06f0;
mem[862] = 144'h0efbf276ff1b019e0dbffd8bfceb0736f59a;
mem[863] = 144'h0ac5f76df50bfab3f1b60cab09a90c78f582;
mem[864] = 144'h00be0310f48f054efd3f099bf592fd260a92;
mem[865] = 144'h05920bdd03740deaf451f81af419fc5df5f5;
mem[866] = 144'hf0e5f027f7b3f3670cfaf18c00660c04f207;
mem[867] = 144'h024bf25701400c15050bffa809dafbadfab2;
mem[868] = 144'hf6f4f0860efd0edeffd10c72f1950d0c0724;
mem[869] = 144'h04200bf10c47084b07470a52fc45f7ba012e;
mem[870] = 144'h0947f16d08b3007d01bd0ba607f2009bf968;
mem[871] = 144'hf164fba7fd590bc6f9befd26fae40b06f901;
mem[872] = 144'hf025f33ffd02fa0cfe10f1d9f598f9a4076a;
mem[873] = 144'h0186f6d10ec9ff9df6a209ec0b79f6160cb4;
mem[874] = 144'h095ff0100274f5e4fa1afcb80da20f700113;
mem[875] = 144'h0f6cfe3b0cf703880e5b0cae0c5402dcf912;
mem[876] = 144'h07a9f170f4d2f120f3870b81018c03d20bbe;
mem[877] = 144'hf5c3f33d073501ac0fee06fbf114ff3ef4d1;
mem[878] = 144'h062df377f183fd4c066a06700cdaf803f588;
mem[879] = 144'h0090fd14051804050a81f81efdb9f00c0022;
mem[880] = 144'h0a9cf4850a4306a206fff19bfe40fa180b60;
mem[881] = 144'h0cdef1d9006707f3f5e40e3202b609acf3b6;
mem[882] = 144'hf22202c8f74af36afd5afe280f1a083affc3;
mem[883] = 144'h02f20732f8380bf605d3f2cffb8702bef279;
mem[884] = 144'hf3b002f0f153009f0b28f08e011e090b0024;
mem[885] = 144'hf4f90a290ee0f3ae098efef50738fb070f58;
mem[886] = 144'hf58cf95dfa0efed809010c0af8fd0213f815;
mem[887] = 144'h0173f18df03bf243f97901cd04ab0a3a05a5;
mem[888] = 144'h0b27f78604e4f9dbf6af0964fd190c73fc71;
mem[889] = 144'h09aef0a50b540b03052bf427fe35f7f8f7e5;
mem[890] = 144'h05820b4805aa09890cb706c4f021f893fb6d;
mem[891] = 144'h0f73fc50f1390399f3b3f683ff790d980b49;
mem[892] = 144'h0e45f281fec60503064defd5f05df7080494;
mem[893] = 144'h0e6af710f1def8c9f30607a7f261faf3f83d;
mem[894] = 144'h0922f6e601e7f850f1c2f0ccff0ff7410bd7;
mem[895] = 144'h08170f0bff47f1ae08d80de7fff3fbd0f328;
mem[896] = 144'h04cf091505abf2680aeaf446f4eefc750db9;
mem[897] = 144'hf0dcf894fae5026c01aa0b7bf5fa0c9ef873;
mem[898] = 144'h0da808d7fb6dfbbff4ed093f04bdf758f75a;
mem[899] = 144'h0653faf0fb36ffaafb4b04510f0d0cdafc61;
mem[900] = 144'hf2bf022ef609f3dd05aef4b8f146ff1a04a0;
mem[901] = 144'h080d0fc403fcf402fcba0c1cf2570628ffd7;
mem[902] = 144'hfa30ff5605d4f023f868f235f2d1fc09006a;
mem[903] = 144'h0bcafffc0c9a01ef0a5c04f700a607de03d5;
mem[904] = 144'h0ae50a98fe7d0d67fb71fe33eff100620375;
mem[905] = 144'hfb6dfa93fd9a0c160e59f360f339f9440ca1;
mem[906] = 144'hf3c9fefc0eeb0c80026106dc0f52056206cf;
mem[907] = 144'h098206a0f9aa00fefc7904850d53f2cff36b;
mem[908] = 144'h095303a904faf9b9f4ff01ff0f6ef7f701df;
mem[909] = 144'hf7160245031404720a56fa320a25fbae0658;
mem[910] = 144'h02410abaf73bfe8ef014fb01f6fbf73b049d;
mem[911] = 144'h0fc609c603c10a5c071df5920a11f39d00da;
mem[912] = 144'h0d9a04a3f92ff2960b64f9dcf55d0a650b7d;
mem[913] = 144'h01580603f008f64bf85bfb28fb13f1e90e72;
mem[914] = 144'hf2cc04ff0d84f7a901440d340393fb62fabc;
mem[915] = 144'hf9b704a0f5bb03650e9c0e5a018df85bf76d;
mem[916] = 144'hf4f0f06400a10d37fe240e76ffff0979f129;
mem[917] = 144'hfa57fbbbfcbdf9970a2f04d5f222ff6af157;
mem[918] = 144'hf8e1fa73fb57082b00d6fa8d020a0b14ffae;
mem[919] = 144'hf959039d0ef9fad6ffb7f4dbf1ed0d190673;
mem[920] = 144'h00ee0ce907b9f1d205cdf1d50d14f80c0338;
mem[921] = 144'hfeda0561ff170d95fd03095c00400c7bf4e8;
mem[922] = 144'h06c30755f1b2f920f57205d4f646f30af035;
mem[923] = 144'hff72fe03071d0e12fae2f75efa07f74a05ff;
mem[924] = 144'hf82afc91f23f04a4f4fb0965f107032bf30b;
mem[925] = 144'h075cffaa0eb305e605bb0aec05ef0c010265;
mem[926] = 144'h08dbf82708baf636f4eff955f7d3f1020059;
mem[927] = 144'h038c04a20023fec5fba6f0190b12f10cf369;
mem[928] = 144'hfbe607e90844f9c2f8e001ec02eafc74fc94;
mem[929] = 144'h0dc90d9d009b0276ff41fecb0553efd6f2bf;
mem[930] = 144'hfa9900e40011fb130ddb00d8ff04fb9c01a4;
mem[931] = 144'hfc89ff61fb3106f3f79cff39089c0e3cff85;
mem[932] = 144'h09aa02df0481fe9affe506dcf6b90c05f634;
mem[933] = 144'hf788001efe25fc0a061c018601090a08f37d;
mem[934] = 144'hf315f249f249006c04bef760f26efb41f20a;
mem[935] = 144'hf1da0e480fb3f57103bb0b82f9a6fe67038c;
mem[936] = 144'hff0cf3a1f34b065e08a60f14fdc30e090c91;
mem[937] = 144'hfe520e6e0a04f4c5f16af9dcfd5a0f940cb7;
mem[938] = 144'hfbf802020d710985f25f005cfb5708c10473;
mem[939] = 144'hf920fc28fdb4ffdaf93f03c2f5600d16fd25;
mem[940] = 144'h0ff00ec0fb34fe1b0462f132f632013803cb;
mem[941] = 144'h0bb8f9180b6003b00eb0fdd0f2c0fc6b0bbb;
mem[942] = 144'h03f7effbf48e064a04f5f6d1052700d20609;
mem[943] = 144'hff59f6fff075fafe078ff4e90a74f7dcf883;
mem[944] = 144'hf9390a1f05230aebfd47fba20f89fe93f501;
mem[945] = 144'hfd6cfc5a0093013bf2a0f31c0593078e0511;
mem[946] = 144'h00bb0a3409a3f7fc04f809b7027df88c07b9;
mem[947] = 144'hfaa4fc17f5d6f47a07d7030f05ac0769062c;
mem[948] = 144'h0ed4fb86fae70cc8f4f9f9ceff3b058307fc;
mem[949] = 144'h068207b9effb04e80d10005afc14fa53feda;
mem[950] = 144'h0dd2fa680d1afde8f57e0a8808700b0fff37;
mem[951] = 144'h02d707bc0d4d0a420554fcccff92065afe26;
mem[952] = 144'hf277f562f4e6ffcffa9ef97b074709920ecf;
mem[953] = 144'h068ff15dfd36f0c9fe96f25c08d1f27405d6;
mem[954] = 144'hf73bf0d1f96a0bf30144f2440f4ef01cf3e2;
mem[955] = 144'hff0203ae078b077603640c9c0beb0f5bf96f;
mem[956] = 144'hfa0d0f59f6b70221f6cbfbd6fde10202f780;
mem[957] = 144'hf2dd00bfffd0fdb8ff2d0bbcf4acf5d3fad8;
mem[958] = 144'h0d1e09190186f0840d490d1a0aaafb0e04ba;
mem[959] = 144'hf7fffc370e10f754f26cf1120c2df6c30c72;
mem[960] = 144'h09d908d6f1df019101bef756fc9f04280df9;
mem[961] = 144'h0eea00e8fbdaf61d0dc207230f35fec9f20d;
mem[962] = 144'hf7e20ec9fb34fc62fca101ff0d25fac9fd2e;
mem[963] = 144'hf412fa6a0ab502a8fc7702dbf680f015f455;
mem[964] = 144'hf64cf0d004bff95306520a7f04edf240f9dc;
mem[965] = 144'hfa62fcb7faae0b160482fd87fbe6f2f3f537;
mem[966] = 144'hf66ff3c6f33b0f24f636f41e0697fd4c0a1c;
mem[967] = 144'hf6010c43f5cd02e8f64309a0055c05980744;
mem[968] = 144'hfc0a0d9c01bf006cf07bf68ef31df3240256;
mem[969] = 144'h09c306aef026f63909d70f1f0d30fb0b0eeb;
mem[970] = 144'h08c30be302d4f60d0aa70242ff67038b08c0;
mem[971] = 144'hfe85f0e6f44207c90851ffddfe3e04e8f5ad;
mem[972] = 144'h09d0fa8d0c08facb010c0523f7bef71b016a;
mem[973] = 144'hf1490ac6f5db0a26091708eb09d0f43708e2;
mem[974] = 144'h055bf181fccbf57afbdd010c08f9047f06da;
mem[975] = 144'hf3840185fcd305a0045ff5cdf2a4f862080a;
mem[976] = 144'h0d32020b0e53025506ce069506b005660ee7;
mem[977] = 144'h0f5ffd1cff0808eef697f353fc24f6fc0ce0;
mem[978] = 144'h015efa09feadfd79f8490807fc09f2c8003e;
mem[979] = 144'hf2c5f34cfc48f63d0b08f7350ab50b300a72;
mem[980] = 144'h08e50f50fb5f0907f68c09daf191f3fb07f8;
mem[981] = 144'h007c0dc1089108e9052909fc0f1d0a77fe8f;
mem[982] = 144'hfdcbf48c07ecfb35f4fb0c32f09df74c051b;
mem[983] = 144'hf975fe6901e60a0dfd2cf5da0fe1fd030f6b;
mem[984] = 144'h00bf0c79fd29fe6df51f03b1f2ae0f89fad3;
mem[985] = 144'hf715f754f2a104550edbf77c05a5f2b2fd0e;
mem[986] = 144'hfe1bfe05f642fccff48ffc13f557f8d50132;
mem[987] = 144'h0da5fb6a0fda0ff4f84afda90b2ffdac0822;
mem[988] = 144'h0766f2d201a9f879fb2ffc580534f6340bf4;
mem[989] = 144'h0d6afb29fea602860829034308cffeb3f5b2;
mem[990] = 144'h0be40375000c04590c800c740125fa530911;
mem[991] = 144'hf9da031ffc4d0e36f50bfa4904820f44f54e;
mem[992] = 144'h09580b7e0efffb7bf89cf7a1f91ff6acf89e;
mem[993] = 144'hf1a9023d0c990573fa3f09f6f9f205ee0eb3;
mem[994] = 144'h08e1097b0e6e04750b17f03cf74bfe71f41e;
mem[995] = 144'h015dfba1f037f201fbd005590b7906050db0;
mem[996] = 144'hf0d8f43a0b36f1c805a20ced0b76fd9c0b43;
mem[997] = 144'hfdacfd7104820639f05304890696fd600394;
mem[998] = 144'hf134fbbc08f6f6460f79f610f63306caf625;
mem[999] = 144'hf74f024dffc3fab102cd0f61042e0d0200de;
mem[1000] = 144'h0edb0f49fa780aa5f92c092208cbf3830bf0;
mem[1001] = 144'hf965f4e1fe4507caf3e0f5cd02b003ec0d57;
mem[1002] = 144'h06ce06bb0392064e0cbb09010e7bfd0a02f7;
mem[1003] = 144'hf07cfe170160ff62fcbe0dbcf4960adefcdc;
mem[1004] = 144'h06f2084f0c330c9effff023d008700640a9a;
mem[1005] = 144'h0d2404d8f168fb68071bfc34f5fafc2400e6;
mem[1006] = 144'h0d33f2fb0bdf04a90edff56f0c930adc0523;
mem[1007] = 144'hf378fdbe02f7f31dfa3e0089065afcd0f50a;
mem[1008] = 144'h04c80182f7a30317f3cc08fe0143f7f80e83;
mem[1009] = 144'hffa3003bf9b6f1e8fbe804090d1c0fe00e60;
mem[1010] = 144'h00b3f920f44109330e3dff41fd8dfe8cf6db;
mem[1011] = 144'hfa29fbf7f9bbf20b06a4f4e9f14901fd0a5c;
mem[1012] = 144'hf3a4019e015ef6c9f3fb0491f143090bf32d;
mem[1013] = 144'h0956f125fe1dff510b74f5acfadbf81af376;
mem[1014] = 144'h0567080cfb11ff22f7c90adc0575f2c50e73;
mem[1015] = 144'h03f703b20b970cc1fc320b5008730b5708c8;
mem[1016] = 144'hfdd005f9f6befef3fd3905490d56008a0e71;
mem[1017] = 144'h0f2507960e96f9cefcd90ab1ffd7f7e0fa43;
mem[1018] = 144'h0f19f21c045c04d3fc7e07830f3e0f77f3d1;
mem[1019] = 144'hf06608d0074afcad0d07f01ff1cbfbc507b7;
mem[1020] = 144'hf261fcd3fb600342ff75f97406eaf7f7febf;
mem[1021] = 144'h0c7007d0018df587f83e048a07370a61fb34;
mem[1022] = 144'hf5cef7aa0b590760f741fccbf8fffc96f2a6;
mem[1023] = 144'hfee70a7903000631fcfcf5230cb30344fb7d;
mem[1024] = 144'h007a0bd4f86105270dba0477fa1e05a10e6a;
mem[1025] = 144'h0466028f07a0f21a02e6f4c5f8ef0d6c0bb8;
mem[1026] = 144'h0dc5f064f23ef8a3fc10f802f8c1f0edf95e;
mem[1027] = 144'h0fc0ff6a0aa90e13fb0d08b603a8facfff79;
mem[1028] = 144'hf5f80ba1058908d8030e041e047f02da0320;
mem[1029] = 144'h0155f50c0decfc54f5cd0fc1f7cb034ef296;
mem[1030] = 144'hf39b0ba8f07f0c4bfbbcf689fe9ff4d40e5d;
mem[1031] = 144'hf12bf7a9fbcbf3b6035c0a3ef81bf75d0f8d;
mem[1032] = 144'h09dd0760088c0722f9b1f6c9f734f3290797;
mem[1033] = 144'h06770f05f94cfd900366f7b90b92fd87f1b6;
mem[1034] = 144'h0b160e05f877f44af364f139f9b60ba5037b;
mem[1035] = 144'hf60efa2c0019f37ef19c057bfae9f8670c38;
mem[1036] = 144'h0559f0120f84fd440dec078ef35b033bf4c2;
mem[1037] = 144'hf329faf60d480ac605da0f580abff990f805;
mem[1038] = 144'h0cccfcb30092057204dd08e003a2f6c5fc0a;
mem[1039] = 144'h06750109f0a9fc4bf6ff0ea00973fc3f0cec;
mem[1040] = 144'h07da07ef03f8f2a401740638fcc9052e0800;
mem[1041] = 144'h0b890f8ffe0901ee0ab2f61df78a050df3d0;
mem[1042] = 144'hf4b3f30006960b00f223f9d4fe2a0459fe65;
mem[1043] = 144'h0723093df8f300a20beaf6ccf899fa920511;
mem[1044] = 144'h0d9b05d7f835064a08b8f3900033ff1b070f;
mem[1045] = 144'h0d50fb590f3f0191f877ff9d0819026cf081;
mem[1046] = 144'hfdc70b3cf07a01e6ff4f059bffa20ceb0cfa;
mem[1047] = 144'hfe22f3f90cbd02d9f081fcf3f6590204045b;
mem[1048] = 144'h0c900db10737fce0fe9405acfe73f2b70d68;
mem[1049] = 144'hfccafbb8fa9d040ff577f2eafb9c00440426;
mem[1050] = 144'hf9c20910fe8706ddf9950216053f0ddbffa7;
mem[1051] = 144'hffa40ee8025cf1b50d870442fb13f3d90312;
mem[1052] = 144'hfd9a0a8e0a360ebcf2260d63f641f200fd68;
mem[1053] = 144'h0c320f9001e90f3c0dd6fda90e3f0ae50696;
mem[1054] = 144'h057209d8079cf15a035bf173fcb803c00586;
mem[1055] = 144'h0db1f9520254f27cf1440069fd01f266f2e8;
mem[1056] = 144'hf17409a4f787094103f00388007902fa0902;
mem[1057] = 144'hf14b0ebafc3e0307ff4df53c0b0e0843018b;
mem[1058] = 144'hfd4bfa840dd007b1f5c10eb80413f1e7f7b0;
mem[1059] = 144'h0221060f08fef4cb07e5f55207dbf25bfe93;
mem[1060] = 144'h0197f11ef3e20d0d028b0d680277f1140232;
mem[1061] = 144'hf472f1d9ffb302e2f5a300480c500ea9f2b8;
mem[1062] = 144'h0a8cf43cfad6f7eff9a6f6eefb390239fc2e;
mem[1063] = 144'hf6a2f81703b004940072f217f7a00003f8b1;
mem[1064] = 144'h0a5d06f30aecf3b5fa96f344f68701d5057b;
mem[1065] = 144'hfc0c04f3070a03e505ac0fa002cff8cbf643;
mem[1066] = 144'h0dff0e5a08890ccd0d8efa21f4cbf985fc05;
mem[1067] = 144'hf1f2fc31f1fdfb68f1a6f976f1c30fd0004b;
mem[1068] = 144'h07e1f9760b8cf9370c180f450e450437059e;
mem[1069] = 144'hf62a034500000609f2e30c02f7100e3b0880;
mem[1070] = 144'h05ea06c003e50fcb08b40f320163fc91f764;
mem[1071] = 144'h0de5f737f2db0a740d980891f584028c0f89;
mem[1072] = 144'hf254ff200899f55bf14ef4e60326fbba0254;
mem[1073] = 144'hf1ccf956071006fa01330b09ffcb00f0081a;
mem[1074] = 144'hf8f8f9c7f37c0a6f026cf6ad011bf56af86c;
mem[1075] = 144'h06f30b2f010204b0fde60739ff9cfea9fd64;
mem[1076] = 144'hf0fffe16f14c037b05e203f70c21f5c3f786;
mem[1077] = 144'h0cd70af4fe1ef1e80145086bfb08f1effd37;
mem[1078] = 144'hf3040b8406fef87906b0f1f5037605b50474;
mem[1079] = 144'hfc64f76c08b0f1e60145038900940e43033d;
mem[1080] = 144'hffaaff3cf4dffc7bf491062ff3590d4e0df6;
mem[1081] = 144'hfa9a05c2f48b02cfffeefe91f1cd0120f0c6;
mem[1082] = 144'h0e1afbee0a0104b2f33cfd63fdb7fcc4f05d;
mem[1083] = 144'hf71ff0660d6a04280856f8e7f7c2fa480475;
mem[1084] = 144'hfa05fd6cf56c0c8e01b7f0d20e61f45afb06;
mem[1085] = 144'h04d5f02006ab00890248f333036cf017030d;
mem[1086] = 144'h04d908250307f984fdd80cccfef1f758f46d;
mem[1087] = 144'hffd9001efa360679fdeef34302e004690b73;
mem[1088] = 144'hf87e0fdcf4870034083bf87df3cf018af07f;
mem[1089] = 144'h0809f0a30338fed90ec8fb730bbcfae5f46c;
mem[1090] = 144'hf81ef2e9fd28f5b1fca1f2effcf5040bff22;
mem[1091] = 144'hf60a09b303cf0f71ffb3085d0deaf718f278;
mem[1092] = 144'h088efb62feecf36408e6fbbbf60905c10f22;
mem[1093] = 144'h06c8081401ed0c1cf66500940deaf771fc2e;
mem[1094] = 144'hfb630874fdfef01aff5b0e73fc9bf9f7f8b4;
mem[1095] = 144'h07a3f82cf3df04e405d003a005ce0e050768;
mem[1096] = 144'hf2d409c3f586ffa2f82c009b0bed00b30c83;
mem[1097] = 144'hfe3efcff04e0f2fb0b70ff96f5550ccaf97a;
mem[1098] = 144'hf969f5370948fb730d7701a3f50807980a61;
mem[1099] = 144'hfd52f51c013709300a950d04fdf900520deb;
end

always @ (posedge clk) begin
	q_a <= mem[addr_a];
end

always @ (posedge clk) begin
	q_b <= mem[addr_b];
end

endmodule